* SPICE NETLIST
***************************************

.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT mimcap_1p0_sin TOP BOT
.ENDS
***************************************
.SUBCKT mimcap_1p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin TOP BOT
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT na20_g5a_cfp_mac D G S B
.ENDS
***************************************
.SUBCKT na20_g5a_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT na29_g5a_cfp_mac D G S B
.ENDS
***************************************
.SUBCKT na29_g5a_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT na6_g5a_nbl_v2_mac D G S B SUB
.ENDS
***************************************
.SUBCKT nch_hv5_5vnw_ac D G S B
.ENDS
***************************************
.SUBCKT nda29_g3a_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT nda45_g3b_nbl_cfp_mac D G BS SUB
.ENDS
***************************************
.SUBCKT ndio_sbd_mac PLUS MINUS
.ENDS
***************************************
.SUBCKT nld12_g5a_cfp_mac D G BS
.ENDS
***************************************
.SUBCKT nld12_g5a_iso_cfp_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld16_g5a_cfp_mac D G BS
.ENDS
***************************************
.SUBCKT nld16_g5a_iso_cfp_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld20_g5a_cfp_mac D G BS
.ENDS
***************************************
.SUBCKT nld20_g5a_iso_cfp_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld24_g5a_cfp_mac D G BS
.ENDS
***************************************
.SUBCKT nld24_g5a_iso_cfp_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld24_g5a_iso_switch_cfp_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld24_g5a_switch_cfp_mac D G BS
.ENDS
***************************************
.SUBCKT nld36_g5b_nbl_cfp_mac D G BS SUB
.ENDS
***************************************
.SUBCKT nld45_g5b_nbl_cfp_mac D G BS SUB
.ENDS
***************************************
.SUBCKT nld5_g5a_iso_switch_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld6_g5a_de_iso_v2_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld6_g5a_de_mac D G BS
.ENDS
***************************************
.SUBCKT nld6_g5a_sa_iso_v2_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld6_g5a_sa_mac D G BS
.ENDS
***************************************
.SUBCKT nld9_g5a_iso_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld9_g5a_mac D G BS
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_5 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_5_mis PLUS MINUS
.ENDS
***************************************
.SUBCKT npddshnnbl10_ga_bgr8_7t C1 C8 B1 B8 E1 E8 SUB
.ENDS
***************************************
.SUBCKT npddshnnbl10_ga_poly_4t C B E SUB
.ENDS
***************************************
.SUBCKT npddshnnbl2_ga_poly_4t C B E SUB
.ENDS
***************************************
.SUBCKT npddshnnbl5_ga_poly_4t C B E SUB
.ENDS
***************************************
.SUBCKT npwshnnbl10_ga_bgr8_7t C1 C8 B1 B8 E1 E8 SUB
.ENDS
***************************************
.SUBCKT npwshnnbl10_ga_poly_4t C B E SUB
.ENDS
***************************************
.SUBCKT npwshnnbl2_ga_poly_4t C B E SUB
.ENDS
***************************************
.SUBCKT npwshnnbl5_ga_poly_4t C B E SUB
.ENDS
***************************************
.SUBCKT pa12_g5a_nbl_slit_v2_mac D G BS SUB
.ENDS
***************************************
.SUBCKT pa12_g5a_nbl_v2_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa16_g5a_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa16_g5a_nbl_slit_cfp_mac D G BS SUB
.ENDS
***************************************
.SUBCKT pa20_g5a_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa20_g5a_nbl_slit_cfp_mac D G BS SUB
.ENDS
***************************************
.SUBCKT pa29_g5a_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa36_g5b_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa45_g5b_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa6_g5a_de_nbl_v2_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa6_g5a_sa_nbl_v2_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa9_g5a_nbl_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa9_g5a_nbl_slit_mac D G BS SUB
.ENDS
***************************************
.SUBCKT pbhvnwshnnbl_esd_dio_shp_gb_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pbshnnbl_dio_shp_ga_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pch5_as_switch_mac D G BS SUB
.ENDS
***************************************
.SUBCKT pddshnnbl_dio_shp_ga_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_12_pdd_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_12_v4_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_16_v3_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_20_pdd_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_20_v3_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_24_v3_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_29_v3_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_6_v3_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_9_v3_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_gb_36_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_gb_45_cit_v3_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT phvnwpsub10_gb_poly C B E
.ENDS
***************************************
.SUBCKT phvnwpsub2_gb_poly C B E
.ENDS
***************************************
.SUBCKT phvnwpsub5_gb_poly C B E
.ENDS
***************************************
.SUBCKT pnddpsub10_ga_poly C B E
.ENDS
***************************************
.SUBCKT pnddpsub2_ga_poly C B E
.ENDS
***************************************
.SUBCKT pnddpsub5_ga_poly C B E
.ENDS
***************************************
.SUBCKT pnddshp5_nbl_ga_4t C B E SUB
.ENDS
***************************************
.SUBCKT rnod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodrpo_pure5v PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodrpo_pure5v_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1rpo_pure5v PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpo1rpo_pure5v_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwod_pure5v PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_pure5v_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwsti_pure5v PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_pure5v_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodrpo_pure5v PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodrpo_pure5v_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1rpo_pure5v PLUS MINUS
.ENDS
***************************************
.SUBCKT rppo1rpo_pure5v_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1rpo_serp PLUS MINUS
.ENDS
***************************************
.SUBCKT rppo1rpo_serp_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppolyhri1k PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyhri1k_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyhri3d3k PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyhri3d3k_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyhri3d3k_serp PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyhri3d3k_serp_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_dio_ga_12_v2_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT sbd_dio_ga_16_v2_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT sbd_dio_ga_24_v2_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT shpnblshn_dio_shp_gb_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT shpshnnbl_esd_dio_shp_ga_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT zd_dio_ga_nbl_v2_4t PLUS MINUS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT tsmc_c018_sealring_corner_1p5m
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT tsmc_c018_seal_ring_edge_1p5m
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_28
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_29
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_30
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_31
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_32
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_CORNER_VIA
** N=6 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT PCORNER
** N=7 EP=0 IP=12 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT HBK183_PAD_LINE_S
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_NMOS_W26_L075_S
** N=5 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=6 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=5 EP=0 IP=12 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_PMOS_W21_L075_S
** N=5 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=5 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=6 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_POSTGR_RES
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_POSTDRV_PDUW0208SCDG_S 1 2 3 4 5 6 7 8
** N=10 EP=8 IP=57 FDC=48
*.SEEDPROM
M0 7 3 2 8 ND L=7.5e-07 W=2.6e-05 $X=5520 $Y=5590 $D=1
M1 2 9 7 8 ND L=7.5e-07 W=2.6e-05 $X=9930 $Y=5590 $D=1
M2 7 9 2 8 ND L=7.5e-07 W=2.6e-05 $X=11900 $Y=5590 $D=1
M3 2 9 7 8 ND L=7.5e-07 W=2.6e-05 $X=16310 $Y=5590 $D=1
M4 7 9 2 8 ND L=7.5e-07 W=2.6e-05 $X=18280 $Y=5590 $D=1
M5 2 9 7 8 ND L=7.5e-07 W=2.6e-05 $X=22690 $Y=5590 $D=1
M6 7 9 2 8 ND L=7.5e-07 W=2.6e-05 $X=24660 $Y=5590 $D=1
M7 2 9 7 8 ND L=7.5e-07 W=2.6e-05 $X=29070 $Y=5590 $D=1
M8 7 9 2 8 ND L=7.5e-07 W=2.6e-05 $X=31040 $Y=5590 $D=1
M9 2 9 7 8 ND L=7.5e-07 W=2.6e-05 $X=35450 $Y=5590 $D=1
M10 7 9 2 8 ND L=7.5e-07 W=2.6e-05 $X=37420 $Y=5590 $D=1
M11 2 9 7 8 ND L=7.5e-07 W=2.6e-05 $X=41830 $Y=5590 $D=1
M12 7 9 2 8 ND L=7.5e-07 W=2.6e-05 $X=43800 $Y=5590 $D=1
M13 2 9 7 8 ND L=7.5e-07 W=2.6e-05 $X=48210 $Y=5590 $D=1
M14 7 9 2 8 ND L=7.5e-07 W=2.6e-05 $X=50180 $Y=5590 $D=1
M15 2 9 7 8 ND L=7.5e-07 W=2.6e-05 $X=54590 $Y=5590 $D=1
M16 7 9 2 8 ND L=7.5e-07 W=2.6e-05 $X=56560 $Y=5590 $D=1
M17 2 9 7 8 ND L=7.5e-07 W=2.6e-05 $X=60970 $Y=5590 $D=1
M18 7 9 2 8 ND L=7.5e-07 W=2.6e-05 $X=62940 $Y=5590 $D=1
M19 2 6 7 8 ND L=7.5e-07 W=2.6e-05 $X=67350 $Y=5590 $D=1
M20 7 6 2 8 ND L=7.5e-07 W=2.6e-05 $X=69320 $Y=5590 $D=1
M21 2 6 7 8 ND L=7.5e-07 W=2.6e-05 $X=73730 $Y=5590 $D=1
M22 7 4 1 1 PD L=7.5e-07 W=2.1e-05 $X=5520 $Y=52340 $D=17
M23 1 4 7 1 PD L=7.5e-07 W=2.1e-05 $X=9930 $Y=52340 $D=17
M24 7 4 1 1 PD L=7.5e-07 W=2.1e-05 $X=11900 $Y=52340 $D=17
M25 1 4 7 1 PD L=7.5e-07 W=2.1e-05 $X=16310 $Y=52340 $D=17
M26 7 10 1 1 PD L=7.5e-07 W=2.1e-05 $X=18280 $Y=52340 $D=17
M27 1 10 7 1 PD L=7.5e-07 W=2.1e-05 $X=22690 $Y=52340 $D=17
M28 7 10 1 1 PD L=7.5e-07 W=2.1e-05 $X=24660 $Y=52340 $D=17
M29 1 10 7 1 PD L=7.5e-07 W=2.1e-05 $X=29070 $Y=52340 $D=17
M30 7 10 1 1 PD L=7.5e-07 W=2.1e-05 $X=31040 $Y=52340 $D=17
M31 1 10 7 1 PD L=7.5e-07 W=2.1e-05 $X=35450 $Y=52340 $D=17
M32 7 10 1 1 PD L=7.5e-07 W=2.1e-05 $X=37420 $Y=52340 $D=17
M33 1 5 7 1 PD L=7.5e-07 W=2.1e-05 $X=41830 $Y=52340 $D=17
M34 7 5 1 1 PD L=7.5e-07 W=2.1e-05 $X=43800 $Y=52340 $D=17
M35 1 5 7 1 PD L=7.5e-07 W=2.1e-05 $X=48210 $Y=52340 $D=17
M36 7 5 1 1 PD L=7.5e-07 W=2.1e-05 $X=50180 $Y=52340 $D=17
M37 1 5 7 1 PD L=7.5e-07 W=2.1e-05 $X=54590 $Y=52340 $D=17
M38 7 5 1 1 PD L=7.5e-07 W=2.1e-05 $X=56560 $Y=52340 $D=17
M39 1 5 7 1 PD L=7.5e-07 W=2.1e-05 $X=60970 $Y=52340 $D=17
M40 7 5 1 1 PD L=7.5e-07 W=2.1e-05 $X=62940 $Y=52340 $D=17
M41 1 5 7 1 PD L=7.5e-07 W=2.1e-05 $X=67350 $Y=52340 $D=17
M42 7 5 1 1 PD L=7.5e-07 W=2.1e-05 $X=69320 $Y=52340 $D=17
M43 1 5 7 1 PD L=7.5e-07 W=2.1e-05 $X=73730 $Y=52340 $D=17
R44 10 1 526.2 $[PR] $X=34295 $Y=44870 $D=52
R45 2 9 526.2 $[PR] $X=49830 $Y=38370 $D=52
D46 8 1 pnwdio_5_iso AREA=2.10858e-09 pj=0.00020828 $X=1690 $Y=49040 $D=112
D47 8 1 pnwdio_iso AREA=2.0976e-11 pj=1.951e-05 $X=47830 $Y=37690 $D=114
.ENDS
***************************************
.SUBCKT HBK183_COMM_N_1
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_NMOS_W2_L06 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 2 1 4 ND L=6e-07 W=2e-06 $X=790 $Y=0 $D=1
.ENDS
***************************************
.SUBCKT HBK183_PMOS_W2_L06_1
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_NMOS_W7_L06 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 2 1 4 ND L=6e-07 W=7e-06 $X=790 $Y=0 $D=1
.ENDS
***************************************
.SUBCKT HBK183_NMOS_W1_L027 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 2 1 4 N L=2.7e-07 W=1e-06 $X=960 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT HBK183_PMOS_W25_L027
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_PMOS_W4_L06
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_PMOS_W5_L06
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_NMOS_W75_L06 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 2 1 4 ND L=6e-07 W=7.5e-06 $X=790 $Y=0 $D=1
.ENDS
***************************************
.SUBCKT HBK183_NMOS_W1_L06 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 2 1 4 ND L=6e-07 W=1e-06 $X=720 $Y=0 $D=1
.ENDS
***************************************
.SUBCKT HBK183_PMOS_W75_L06
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_NMOS_W5_L06 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 2 1 4 ND L=6e-07 W=5e-06 $X=790 $Y=0 $D=1
.ENDS
***************************************
.SUBCKT HBK183_PMOS_W3_L06_1
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_NMOS_W6_L06 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 2 1 4 ND L=6e-07 W=6e-06 $X=790 $Y=0 $D=1
.ENDS
***************************************
.SUBCKT HBK183_PMOS_W2_L06
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_POC_MOS 1 2 3
** N=3 EP=3 IP=4 FDC=1
X0 1 1 2 3 HBK183_NMOS_W2_L06 $T=0 730 0 0 $X=-450 $Y=-30
.ENDS
***************************************
.SUBCKT HBK183_PMOS_W5_L05
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_NMOS_W5_L056_1 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 ND L=6e-07 W=5e-06 $X=790 $Y=0 $D=1
.ENDS
***************************************
.SUBCKT HBK183_PREDRV 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
** N=43 EP=20 IP=329 FDC=84
*.SEEDPROM
M0 3 40 13 20 N L=2.7e-07 W=2e-06 $X=57065 $Y=24440 $D=0
M1 5 25 3 20 ND L=6e-07 W=5e-06 $X=12720 $Y=17440 $D=1
M2 14 3 3 20 ND L=6e-07 W=2e-06 $X=60170 $Y=24440 $D=1
M3 40 39 3 20 ND L=6e-07 W=2e-06 $X=63250 $Y=24440 $D=1
M4 3 15 39 20 ND L=6e-07 W=5.5e-06 $X=64050 $Y=17440 $D=1
M5 2 4 23 2 P L=2.7e-07 W=2.5e-06 $X=5510 $Y=31240 $D=16
M6 31 7 2 2 P L=2.7e-07 W=2.5e-06 $X=26600 $Y=31240 $D=16
M7 2 10 36 2 P L=2.7e-07 W=2.5e-06 $X=40480 $Y=31240 $D=16
M8 38 11 2 2 P L=2.7e-07 W=2.5e-06 $X=44640 $Y=31240 $D=16
M9 13 40 2 2 P L=2.7e-07 W=2.5e-06 $X=55455 $Y=31240 $D=16
M10 2 40 13 2 P L=2.7e-07 W=2.5e-06 $X=57065 $Y=31240 $D=16
M11 41 16 2 2 P L=2.7e-07 W=2.5e-06 $X=67590 $Y=31240 $D=16
M12 22 21 1 1 PD L=6e-07 W=1e-06 $X=2080 $Y=8100 $D=17
M13 1 24 21 1 PD L=6e-07 W=2e-06 $X=4540 $Y=7100 $D=17
M14 24 21 1 1 PD L=6e-07 W=2e-06 $X=6140 $Y=7100 $D=17
M15 27 24 1 1 PD L=6e-07 W=4e-06 $X=6940 $Y=1600 $D=17
M16 25 26 1 1 PD L=6e-07 W=5e-06 $X=9520 $Y=4100 $D=17
M17 1 22 25 1 PD L=6e-07 W=5e-06 $X=11120 $Y=4100 $D=17
M18 5 25 1 1 PD L=6e-07 W=5e-06 $X=12720 $Y=4100 $D=17
M19 6 28 1 1 PD L=6e-07 W=7.5e-06 $X=15680 $Y=1600 $D=17
M20 1 28 6 1 PD L=6e-07 W=7.5e-06 $X=17280 $Y=1600 $D=17
M21 43 27 1 1 PD L=6e-07 W=3e-06 $X=18880 $Y=6100 $D=17
M22 28 33 43 1 PD L=6e-07 W=3e-06 $X=20480 $Y=6100 $D=17
M23 1 29 26 1 PD L=6e-07 W=5e-06 $X=23060 $Y=1600 $D=17
M24 29 30 1 1 PD L=6e-07 W=4e-06 $X=24660 $Y=1600 $D=17
M25 1 32 30 1 PD L=6e-07 W=2e-06 $X=25640 $Y=7100 $D=17
M26 32 30 1 1 PD L=6e-07 W=2e-06 $X=27240 $Y=7100 $D=17
M27 33 32 1 1 PD L=6e-07 W=4e-06 $X=29580 $Y=1600 $D=17
M28 8 34 6 1 PD L=6e-07 W=7.5e-06 $X=32590 $Y=1600 $D=17
M29 1 35 8 1 PD L=6e-07 W=5e-06 $X=34190 $Y=1600 $D=17
M30 5 34 9 1 PD L=6e-07 W=5e-06 $X=36770 $Y=4100 $D=17
M31 1 34 35 1 PD L=6e-07 W=2e-06 $X=39510 $Y=6390 $D=17
M32 34 35 1 1 PD L=6e-07 W=2e-06 $X=41110 $Y=6390 $D=17
M33 1 12 37 1 PD L=6e-07 W=2e-06 $X=43680 $Y=6390 $D=17
M34 12 37 1 1 PD L=6e-07 W=2e-06 $X=45280 $Y=6390 $D=17
M35 40 39 2 2 PD L=6e-07 W=2e-06 $X=60050 $Y=31240 $D=17
M36 2 39 40 2 PD L=6e-07 W=2e-06 $X=61650 $Y=31240 $D=17
M37 40 39 2 2 PD L=6e-07 W=2e-06 $X=63250 $Y=31240 $D=17
M38 1 15 39 1 PD L=6e-07 W=2e-06 $X=64050 $Y=1600 $D=17
M39 1 14 17 1 PD L=6e-07 W=2e-06 $X=66630 $Y=2370 $D=17
M40 14 17 1 1 PD L=6e-07 W=2e-06 $X=68230 $Y=2370 $D=17
M41 18 1 1 1 PD L=5e-07 W=5e-06 $X=71480 $Y=1600 $D=17
M42 1 1 18 1 PD L=5e-07 W=5e-06 $X=73080 $Y=1600 $D=17
M43 18 1 1 1 PD L=5e-07 W=5e-06 $X=74680 $Y=1600 $D=17
M44 1 1 18 1 PD L=5e-07 W=5e-06 $X=76280 $Y=1600 $D=17
R45 18 19 554.264 $[PR] $X=73740 $Y=31490 $D=52
D46 20 2 pnwdio_5_iso AREA=3.44535e-11 pj=2.368e-05 $X=58810 $Y=29040 $D=112
X56 22 21 3 20 HBK183_NMOS_W2_L06 $T=3470 17440 1 180 $X=840 $Y=16680
X57 29 30 3 20 HBK183_NMOS_W2_L06 $T=22270 24440 0 0 $X=21820 $Y=23680
X60 21 23 3 20 HBK183_NMOS_W7_L06 $T=3750 17440 0 0 $X=3300 $Y=16680
X61 3 4 24 20 HBK183_NMOS_W7_L06 $T=5350 17440 0 0 $X=4900 $Y=16680
X62 3 7 30 20 HBK183_NMOS_W7_L06 $T=27030 17440 1 180 $X=24400 $Y=16680
X63 32 31 3 20 HBK183_NMOS_W7_L06 $T=28630 17440 1 180 $X=26000 $Y=16680
X64 35 36 3 20 HBK183_NMOS_W7_L06 $T=38720 17440 0 0 $X=38270 $Y=16680
X65 3 10 34 20 HBK183_NMOS_W7_L06 $T=40320 17440 0 0 $X=39870 $Y=16680
X66 3 11 37 20 HBK183_NMOS_W7_L06 $T=45070 17440 1 180 $X=42440 $Y=16680
X67 12 38 3 20 HBK183_NMOS_W7_L06 $T=46670 17440 1 180 $X=44040 $Y=16680
X68 3 16 17 20 HBK183_NMOS_W7_L06 $T=68020 17440 1 180 $X=65390 $Y=16680
X69 14 41 3 20 HBK183_NMOS_W7_L06 $T=69620 17440 1 180 $X=66990 $Y=16680
X70 3 4 23 20 HBK183_NMOS_W1_L027 $T=6740 26440 0 180 $X=4290 $Y=24680
X71 3 7 31 20 HBK183_NMOS_W1_L027 $T=25640 26440 1 0 $X=25380 $Y=24680
X72 3 10 36 20 HBK183_NMOS_W1_L027 $T=41710 26440 0 180 $X=39260 $Y=24680
X73 3 11 38 20 HBK183_NMOS_W1_L027 $T=43680 26440 1 0 $X=43420 $Y=24680
X74 3 16 41 20 HBK183_NMOS_W1_L027 $T=66630 26440 1 0 $X=66370 $Y=24680
X97 42 26 25 20 HBK183_NMOS_W75_L06 $T=10910 17440 1 180 $X=8280 $Y=16680
X98 3 22 42 20 HBK183_NMOS_W75_L06 $T=12510 17440 1 180 $X=9880 $Y=16680
X99 3 24 27 20 HBK183_NMOS_W1_L06 $T=11940 25440 0 0 $X=11490 $Y=24720
X100 27 24 3 20 HBK183_NMOS_W1_L06 $T=13400 25440 0 0 $X=12950 $Y=24720
X101 33 32 3 20 HBK183_NMOS_W1_L06 $T=30970 17440 1 180 $X=28480 $Y=16720
X105 3 28 6 20 HBK183_NMOS_W5_L06 $T=14890 17440 0 0 $X=14440 $Y=16680
X106 6 28 3 20 HBK183_NMOS_W5_L06 $T=16490 17440 0 0 $X=16040 $Y=16680
X107 26 29 3 20 HBK183_NMOS_W5_L06 $T=22270 17440 0 0 $X=21820 $Y=16680
X108 6 35 8 20 HBK183_NMOS_W5_L06 $T=31800 17440 0 0 $X=31350 $Y=16680
X109 5 35 9 20 HBK183_NMOS_W5_L06 $T=34380 17440 0 0 $X=33930 $Y=16680
X110 9 34 3 20 HBK183_NMOS_W5_L06 $T=35980 17440 0 0 $X=35530 $Y=16680
X113 3 27 28 20 HBK183_NMOS_W6_L06 $T=18090 17440 0 0 $X=17640 $Y=16680
X114 3 33 28 20 HBK183_NMOS_W6_L06 $T=21870 17440 1 180 $X=19240 $Y=16680
X127 3 24 20 HBK183_POC_MOS $T=31110 23710 1 180 $X=28480 $Y=23680
X128 3 35 20 HBK183_POC_MOS $T=35980 23710 0 0 $X=35530 $Y=23680
X129 3 12 20 HBK183_POC_MOS $T=51540 23710 1 180 $X=48910 $Y=23680
X134 3 18 3 20 HBK183_NMOS_W5_L056_1 $T=70640 21440 0 0 $X=70190 $Y=20680
X135 18 3 3 20 HBK183_NMOS_W5_L056_1 $T=72240 21440 0 0 $X=71790 $Y=20680
X136 3 18 3 20 HBK183_NMOS_W5_L056_1 $T=73840 21440 0 0 $X=73390 $Y=20680
X137 18 3 3 20 HBK183_NMOS_W5_L056_1 $T=75440 21440 0 0 $X=74990 $Y=20680
.ENDS
***************************************
.SUBCKT HBK183_M3456
** N=6 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT PAD70LU_TRL
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_PMOS_W45_L06
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_PMOS_W15_L06_1
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_NMOS_W3_L06 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 2 1 4 ND L=6e-07 W=3e-06 $X=790 $Y=0 $D=1
.ENDS
***************************************
.SUBCKT HBK183_SCH_CELL 1 2 3 4 5
** N=8 EP=5 IP=48 FDC=5
X0 7 4 3 1 HBK183_NMOS_W2_L06 $T=10580 17910 0 0 $X=10130 $Y=17150
X8 1 2 6 1 HBK183_NMOS_W3_L06 $T=3490 16910 1 180 $X=860 $Y=16150
X9 6 2 1 1 HBK183_NMOS_W3_L06 $T=5090 16910 1 180 $X=2460 $Y=16150
X10 7 5 6 1 HBK183_NMOS_W3_L06 $T=6690 16910 1 180 $X=4060 $Y=16150
X11 4 5 7 1 HBK183_NMOS_W3_L06 $T=8290 16910 1 180 $X=5660 $Y=16150
.ENDS
***************************************
.SUBCKT HBK183_PUCELL_N 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 1 2 4 ND L=6.6e-06 W=6e-07 $X=1450 $Y=5060 $D=1
.ENDS
***************************************
.SUBCKT PFILLER0005
** N=6 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_71
** N=4 EP=0 IP=12 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT PDDW0208CDG VDDPST VDD VSS VSSPST PAD OEN I DS IE C PE 13
** N=25 EP=12 IP=86 FDC=145
*.SEEDPROM
M0 VDDPST 17 18 VDDPST PD L=6e-07 W=4.5e-06 $X=50150 $Y=82610 $D=17
M1 15 14 VDDPST VDDPST PD L=6e-07 W=1.5e-06 $X=50150 $Y=88610 $D=17
M2 18 17 VDDPST VDDPST PD L=6e-07 W=4.5e-06 $X=51750 $Y=82610 $D=17
M3 VDDPST 14 15 VDDPST PD L=6e-07 W=1.5e-06 $X=51750 $Y=88610 $D=17
M4 15 17 18 VDDPST PD L=6e-07 W=4.5e-06 $X=53350 $Y=82610 $D=17
M5 18 17 15 VDDPST PD L=6e-07 W=4.5e-06 $X=54950 $Y=82610 $D=17
M6 VDDPST VDDPST VDDPST VDDPST PD L=6e-07 W=5e-06 $X=59420 $Y=82610 $D=17
X7 VDDPST VSSPST 19 20 21 22 PAD 13 HBK183_POSTDRV_PDUW0208SCDG_S $T=0 0 0 0 $X=-600 $Y=0
X8 VSS VSS VSS 13 HBK183_NMOS_W2_L06 $T=58630 99500 0 0 $X=58180 $Y=98740
X10 VDDPST VDD VSS OEN 19 20 I 21 22 DS IE 14 C 24 15 PE 23 17 PAD 13 HBK183_PREDRV $T=0 81010 0 0 $X=-600 $Y=80290
X18 VSS 14 16 13 HBK183_NMOS_W3_L06 $T=51540 98500 1 180 $X=48910 $Y=97740
X19 16 14 VSS 13 HBK183_NMOS_W3_L06 $T=53140 98500 1 180 $X=50510 $Y=97740
X20 25 17 16 13 HBK183_NMOS_W3_L06 $T=54740 98500 1 180 $X=52110 $Y=97740
X21 15 17 25 13 HBK183_NMOS_W3_L06 $T=56340 98500 1 180 $X=53710 $Y=97740
X22 24 17 VSS 13 HBK183_PUCELL_N $T=69190 93910 0 0 $X=69130 $Y=93910
.ENDS
***************************************
.SUBCKT HBK183_POSTDRV_GR_VDD2DYN_S
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT HBK183_PREDRV_GR_VDD2DYN_S
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT HBK183_DYNVDD2_LINE_VDD_S
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_DYNVDD2_LINE_VDDPST
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_PAD_LINE_VDD2DYN_S
** N=4 EP=0 IP=54 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_NMOS_W26_L06_DYN_VDD2_S
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_19
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_20
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_RES_8X024_DYN_S
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_NMOS_5X2_S
** N=5 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_NMOS_W15_L6D3_DYN_2
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT PVDD2CDG VDDPST VSSPST VSS 6
** N=10 EP=4 IP=96 FDC=60
*.SEEDPROM
M0 VDDPST 9 VSSPST 6 ND L=6e-07 W=2.6e-05 $X=4130 $Y=5590 $D=1
M1 VDDPST 7 VSS 6 ND L=6e-07 W=2.6e-05 $X=4130 $Y=85680 $D=1
M2 VSSPST 9 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=8390 $Y=5590 $D=1
M3 VSS 7 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=8390 $Y=85680 $D=1
M4 VDDPST 9 VSSPST 6 ND L=6e-07 W=2.6e-05 $X=10210 $Y=5590 $D=1
M5 VDDPST 7 VSS 6 ND L=6e-07 W=2.6e-05 $X=10210 $Y=85680 $D=1
M6 VSSPST 9 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=14470 $Y=5590 $D=1
M7 VSS 7 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=14470 $Y=85680 $D=1
M8 VDDPST 9 VSSPST 6 ND L=6e-07 W=2.6e-05 $X=16290 $Y=5590 $D=1
M9 VDDPST 7 VSS 6 ND L=6e-07 W=2.6e-05 $X=16290 $Y=85680 $D=1
M10 VSSPST 8 7 VSSPST ND L=1e-06 W=1e-06 $X=20320 $Y=75070 $D=1
M11 VSSPST 9 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=20550 $Y=5590 $D=1
M12 VSS 7 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=20550 $Y=85680 $D=1
M13 VDDPST 9 VSSPST 6 ND L=6e-07 W=2.6e-05 $X=22370 $Y=5590 $D=1
M14 VDDPST 7 VSS 6 ND L=6e-07 W=2.6e-05 $X=22370 $Y=85680 $D=1
M15 VSSPST 8 VSSPST VSSPST ND L=6.3e-06 W=1.683e-05 $X=22740 $Y=47370 $D=1
M16 VSSPST 8 VSSPST VSSPST ND L=6.3e-06 W=1.683e-05 $X=22740 $Y=54970 $D=1
M17 VSSPST 8 VSSPST VSSPST ND L=6.3e-06 W=1.683e-05 $X=22740 $Y=62570 $D=1
M18 VSSPST 8 VSSPST VSSPST ND L=6.3e-06 W=1.683e-05 $X=22740 $Y=70170 $D=1
M19 VSSPST 9 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=26630 $Y=5590 $D=1
M20 VSS 7 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=26630 $Y=85680 $D=1
M21 VDDPST 9 VSSPST 6 ND L=6e-07 W=2.6e-05 $X=28450 $Y=5590 $D=1
M22 VDDPST 7 VSS 6 ND L=6e-07 W=2.6e-05 $X=28450 $Y=85680 $D=1
M23 VSSPST 9 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=32710 $Y=5590 $D=1
M24 VSS 7 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=32710 $Y=85680 $D=1
M25 VDDPST 9 VSSPST 6 ND L=6e-07 W=2.6e-05 $X=34530 $Y=5590 $D=1
M26 VDDPST 7 VSS 6 ND L=6e-07 W=2.6e-05 $X=34530 $Y=85680 $D=1
M27 VSSPST 9 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=38790 $Y=5590 $D=1
M28 VSS 7 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=38790 $Y=85680 $D=1
M29 VSSPST 8 VSSPST VSSPST ND L=6.3e-06 W=1.683e-05 $X=40430 $Y=47370 $D=1
M30 VSSPST 8 VSSPST VSSPST ND L=6.3e-06 W=1.683e-05 $X=40430 $Y=54970 $D=1
M31 VSSPST 8 VSSPST VSSPST ND L=6.3e-06 W=1.683e-05 $X=40430 $Y=62570 $D=1
M32 VSSPST 8 VSSPST VSSPST ND L=6.3e-06 W=1.683e-05 $X=40430 $Y=70170 $D=1
M33 VDDPST 9 VSSPST 6 ND L=6e-07 W=2.6e-05 $X=40610 $Y=5590 $D=1
M34 VDDPST 7 VSS 6 ND L=6e-07 W=2.6e-05 $X=40610 $Y=85680 $D=1
M35 VSSPST 9 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=44870 $Y=5590 $D=1
M36 VSS 7 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=44870 $Y=85680 $D=1
M37 VDDPST 9 VSSPST 6 ND L=6e-07 W=2.6e-05 $X=46690 $Y=5590 $D=1
M38 VDDPST 7 VSS 6 ND L=6e-07 W=2.6e-05 $X=46690 $Y=85680 $D=1
M39 VSSPST 9 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=50950 $Y=5590 $D=1
M40 VSS 7 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=50950 $Y=85680 $D=1
M41 VDDPST 9 VSSPST 6 ND L=6e-07 W=2.6e-05 $X=52770 $Y=5590 $D=1
M42 VDDPST 7 VSS 6 ND L=6e-07 W=2.6e-05 $X=52770 $Y=85680 $D=1
M43 VSSPST 9 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=57030 $Y=5590 $D=1
M44 VSS 7 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=57030 $Y=85680 $D=1
M45 9 8 VSSPST VSSPST ND L=1e-06 W=1e-06 $X=58680 $Y=46890 $D=1
M46 VDDPST 9 VSSPST 6 ND L=6e-07 W=2.6e-05 $X=58850 $Y=5590 $D=1
M47 VDDPST 7 VSS 6 ND L=6e-07 W=2.6e-05 $X=58850 $Y=85680 $D=1
M48 VSSPST 9 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=63110 $Y=5590 $D=1
M49 VSS 7 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=63110 $Y=85680 $D=1
M50 VDDPST 9 VSSPST 6 ND L=6e-07 W=2.6e-05 $X=64930 $Y=5590 $D=1
M51 VDDPST 7 VSS 6 ND L=6e-07 W=2.6e-05 $X=64930 $Y=85680 $D=1
M52 VSSPST 9 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=69190 $Y=5590 $D=1
M53 VSS 7 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=69190 $Y=85680 $D=1
M54 VDDPST 9 VSSPST 6 ND L=6e-07 W=2.6e-05 $X=71010 $Y=5590 $D=1
M55 VDDPST 7 VSS 6 ND L=6e-07 W=2.6e-05 $X=71010 $Y=85680 $D=1
M56 VSSPST 9 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=75270 $Y=5590 $D=1
M57 VSS 7 VDDPST 6 ND L=6e-07 W=2.6e-05 $X=75270 $Y=85680 $D=1
R58 10 8 820578 $[PR] $X=6900 $Y=45810 $D=52
R59 10 VDDPST 805174 $[PR] $X=59280 $Y=50110 $D=52
.ENDS
***************************************
.SUBCKT HBK183_PREDRV_GR_VSS3DYN_S
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT HBK183_DYNVDD2_LINE_VSS_S
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_DYNVDD2_LINE_VSSPST_S
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_57
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_58
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_PAD_LINE_VSS3DYN_S
** N=2 EP=0 IP=32 FDC=0
.ENDS
***************************************
.SUBCKT PVSS3CDG VDDPST VSS
** N=8 EP=2 IP=92 FDC=60
*.SEEDPROM
M0 VDDPST 7 VSS VSS ND L=6e-07 W=2.6e-05 $X=4130 $Y=5590 $D=1
M1 VDDPST 5 VSS VSS ND L=6e-07 W=2.6e-05 $X=4130 $Y=85680 $D=1
M2 VSS 7 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=8390 $Y=5590 $D=1
M3 VSS 5 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=8390 $Y=85680 $D=1
M4 VDDPST 7 VSS VSS ND L=6e-07 W=2.6e-05 $X=10210 $Y=5590 $D=1
M5 VDDPST 5 VSS VSS ND L=6e-07 W=2.6e-05 $X=10210 $Y=85680 $D=1
M6 VSS 7 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=14470 $Y=5590 $D=1
M7 VSS 5 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=14470 $Y=85680 $D=1
M8 VDDPST 7 VSS VSS ND L=6e-07 W=2.6e-05 $X=16290 $Y=5590 $D=1
M9 VDDPST 5 VSS VSS ND L=6e-07 W=2.6e-05 $X=16290 $Y=85680 $D=1
M10 VSS 6 5 VSS ND L=1e-06 W=1e-06 $X=20320 $Y=75070 $D=1
M11 VSS 7 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=20550 $Y=5590 $D=1
M12 VSS 5 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=20550 $Y=85680 $D=1
M13 VDDPST 7 VSS VSS ND L=6e-07 W=2.6e-05 $X=22370 $Y=5590 $D=1
M14 VDDPST 5 VSS VSS ND L=6e-07 W=2.6e-05 $X=22370 $Y=85680 $D=1
M15 VSS 6 VSS VSS ND L=6.3e-06 W=1.683e-05 $X=22740 $Y=47370 $D=1
M16 VSS 6 VSS VSS ND L=6.3e-06 W=1.683e-05 $X=22740 $Y=54970 $D=1
M17 VSS 6 VSS VSS ND L=6.3e-06 W=1.683e-05 $X=22740 $Y=62570 $D=1
M18 VSS 6 VSS VSS ND L=6.3e-06 W=1.683e-05 $X=22740 $Y=70170 $D=1
M19 VSS 7 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=26630 $Y=5590 $D=1
M20 VSS 5 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=26630 $Y=85680 $D=1
M21 VDDPST 7 VSS VSS ND L=6e-07 W=2.6e-05 $X=28450 $Y=5590 $D=1
M22 VDDPST 5 VSS VSS ND L=6e-07 W=2.6e-05 $X=28450 $Y=85680 $D=1
M23 VSS 7 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=32710 $Y=5590 $D=1
M24 VSS 5 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=32710 $Y=85680 $D=1
M25 VDDPST 7 VSS VSS ND L=6e-07 W=2.6e-05 $X=34530 $Y=5590 $D=1
M26 VDDPST 5 VSS VSS ND L=6e-07 W=2.6e-05 $X=34530 $Y=85680 $D=1
M27 VSS 7 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=38790 $Y=5590 $D=1
M28 VSS 5 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=38790 $Y=85680 $D=1
M29 VSS 6 VSS VSS ND L=6.3e-06 W=1.683e-05 $X=40430 $Y=47370 $D=1
M30 VSS 6 VSS VSS ND L=6.3e-06 W=1.683e-05 $X=40430 $Y=54970 $D=1
M31 VSS 6 VSS VSS ND L=6.3e-06 W=1.683e-05 $X=40430 $Y=62570 $D=1
M32 VSS 6 VSS VSS ND L=6.3e-06 W=1.683e-05 $X=40430 $Y=70170 $D=1
M33 VDDPST 7 VSS VSS ND L=6e-07 W=2.6e-05 $X=40610 $Y=5590 $D=1
M34 VDDPST 5 VSS VSS ND L=6e-07 W=2.6e-05 $X=40610 $Y=85680 $D=1
M35 VSS 7 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=44870 $Y=5590 $D=1
M36 VSS 5 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=44870 $Y=85680 $D=1
M37 VDDPST 7 VSS VSS ND L=6e-07 W=2.6e-05 $X=46690 $Y=5590 $D=1
M38 VDDPST 5 VSS VSS ND L=6e-07 W=2.6e-05 $X=46690 $Y=85680 $D=1
M39 VSS 7 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=50950 $Y=5590 $D=1
M40 VSS 5 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=50950 $Y=85680 $D=1
M41 VDDPST 7 VSS VSS ND L=6e-07 W=2.6e-05 $X=52770 $Y=5590 $D=1
M42 VDDPST 5 VSS VSS ND L=6e-07 W=2.6e-05 $X=52770 $Y=85680 $D=1
M43 VSS 7 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=57030 $Y=5590 $D=1
M44 VSS 5 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=57030 $Y=85680 $D=1
M45 7 6 VSS VSS ND L=1e-06 W=1e-06 $X=58680 $Y=46890 $D=1
M46 VDDPST 7 VSS VSS ND L=6e-07 W=2.6e-05 $X=58850 $Y=5590 $D=1
M47 VDDPST 5 VSS VSS ND L=6e-07 W=2.6e-05 $X=58850 $Y=85680 $D=1
M48 VSS 7 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=63110 $Y=5590 $D=1
M49 VSS 5 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=63110 $Y=85680 $D=1
M50 VDDPST 7 VSS VSS ND L=6e-07 W=2.6e-05 $X=64930 $Y=5590 $D=1
M51 VDDPST 5 VSS VSS ND L=6e-07 W=2.6e-05 $X=64930 $Y=85680 $D=1
M52 VSS 7 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=69190 $Y=5590 $D=1
M53 VSS 5 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=69190 $Y=85680 $D=1
M54 VDDPST 7 VSS VSS ND L=6e-07 W=2.6e-05 $X=71010 $Y=5590 $D=1
M55 VDDPST 5 VSS VSS ND L=6e-07 W=2.6e-05 $X=71010 $Y=85680 $D=1
M56 VSS 7 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=75270 $Y=5590 $D=1
M57 VSS 5 VDDPST VSS ND L=6e-07 W=2.6e-05 $X=75270 $Y=85680 $D=1
R58 8 6 820578 $[PR] $X=6900 $Y=45810 $D=52
R59 8 VDDPST 805174 $[PR] $X=59280 $Y=50110 $D=52
.ENDS
***************************************
.SUBCKT __$$VIA34_520_520_58_21
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_85 2 3 4 5 6 7 8 9 10
** N=21 EP=9 IP=156 FDC=410
*.SEEDPROM
M0 4 20 21 4 PD L=6e-07 W=4.5e-06 $X=180150 $Y=82610 $D=17
M1 17 16 4 4 PD L=6e-07 W=1.5e-06 $X=180150 $Y=88610 $D=17
M2 21 20 4 4 PD L=6e-07 W=4.5e-06 $X=181750 $Y=82610 $D=17
M3 4 16 17 4 PD L=6e-07 W=1.5e-06 $X=181750 $Y=88610 $D=17
M4 17 20 21 4 PD L=6e-07 W=4.5e-06 $X=183350 $Y=82610 $D=17
M5 21 20 17 4 PD L=6e-07 W=4.5e-06 $X=184950 $Y=82610 $D=17
M6 21 17 5 4 PD L=6e-07 W=5e-06 $X=189420 $Y=82610 $D=17
X36 4 5 12 13 14 15 2 5 HBK183_POSTDRV_PDUW0208SCDG_S $T=130000 0 0 0 $X=129400 $Y=0
X37 4 6 5 7 12 13 8 14 15 8 7 16 10 19 17 7 18 20 2 5 HBK183_PREDRV $T=130000 81010 0 0 $X=129400 $Y=80290
X43 5 16 4 17 20 HBK183_SCH_CELL $T=178050 81590 0 0 $X=176245 $Y=81220
X44 19 20 5 5 HBK183_PUCELL_N $T=199190 93910 0 0 $X=199130 $Y=93910
X56 4 6 5 5 3 7 8 8 7 9 7 5 PDDW0208CDG $T=210030 0 0 0 $X=209430 $Y=0
X57 4 5 5 5 PVDD2CDG $T=290065 0 0 0 $X=289465 $Y=0
X58 4 5 PVSS3CDG $T=370100 0 0 0 $X=369500 $Y=0
.ENDS
***************************************
.SUBCKT TAPCELLBWP7T
** N=2 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT FILL1BWP7T
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_49
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT DCAPBWP7T VDD VSS
** N=4 EP=2 IP=0 FDC=2
*.SEEDPROM
M0 3 4 VSS VSS N L=1.8e-07 W=1e-06 $X=800 $Y=345 $D=0
M1 4 3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=680 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT DCAP8BWP7T VSS VDD
** N=4 EP=2 IP=0 FDC=6
*.SEEDPROM
M0 VSS 4 VSS VSS N L=9.9e-07 W=9.45e-07 $X=620 $Y=345 $D=0
M1 VSS 4 VSS VSS N L=9.9e-07 W=9.45e-07 $X=2150 $Y=345 $D=0
M2 3 4 VSS VSS N L=1.8e-07 W=9.45e-07 $X=3680 $Y=345 $D=0
M3 VDD 3 VDD VDD P L=9.9e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M4 VDD 3 VDD VDD P L=9.9e-07 W=1.235e-06 $X=2150 $Y=2340 $D=16
M5 4 3 VDD VDD P L=1.8e-07 W=1.235e-06 $X=3680 $Y=2340 $D=16
.ENDS
***************************************
.SUBCKT DCAP4BWP7T VSS VDD
** N=4 EP=2 IP=0 FDC=4
*.SEEDPROM
M0 VSS 4 VSS VSS N L=2.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 3 4 VSS VSS N L=1.8e-07 W=1e-06 $X=1440 $Y=345 $D=0
M2 VDD 3 VDD VDD P L=2.8e-07 W=1.17e-06 $X=620 $Y=2405 $D=16
M3 4 3 VDD VDD P L=1.8e-07 W=1.17e-06 $X=1440 $Y=2405 $D=16
.ENDS
***************************************
.SUBCKT ICV_40 1 2
** N=2 EP=2 IP=4 FDC=10
*.SEEDPROM
X0 1 2 DCAP8BWP7T $T=0 0 0 0 $X=-290 $Y=-235
X1 1 2 DCAP4BWP7T $T=4480 0 0 0 $X=4190 $Y=-235
.ENDS
***************************************
.SUBCKT NR2D1BWP7T A2 VDD ZN A1 VSS
** N=6 EP=5 IP=0 FDC=4
*.SEEDPROM
M0 ZN A2 VSS VSS N L=1.8e-07 W=1e-06 $X=660 $Y=345 $D=0
M1 VSS A1 ZN VSS N L=1.8e-07 W=1e-06 $X=1420 $Y=345 $D=0
M2 6 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M3 ZN A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=1260 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT DCAP64BWP7T VDD VSS
** N=4 EP=2 IP=0 FDC=48
*.SEEDPROM
M0 VSS 3 4 VSS N L=1.8e-07 W=9.4e-07 $X=620 $Y=405 $D=0
M1 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=1340 $Y=405 $D=0
M2 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=2870 $Y=405 $D=0
M3 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=4400 $Y=405 $D=0
M4 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=5930 $Y=405 $D=0
M5 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=7460 $Y=405 $D=0
M6 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=8990 $Y=405 $D=0
M7 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=10520 $Y=405 $D=0
M8 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=12050 $Y=405 $D=0
M9 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=13580 $Y=405 $D=0
M10 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=15110 $Y=405 $D=0
M11 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=16640 $Y=405 $D=0
M12 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=18170 $Y=405 $D=0
M13 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=19700 $Y=405 $D=0
M14 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=21230 $Y=405 $D=0
M15 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=22760 $Y=405 $D=0
M16 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=24290 $Y=405 $D=0
M17 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=25820 $Y=405 $D=0
M18 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=27350 $Y=405 $D=0
M19 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=28880 $Y=405 $D=0
M20 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=30410 $Y=405 $D=0
M21 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=31940 $Y=405 $D=0
M22 VSS 3 VSS VSS N L=9.9e-07 W=9.4e-07 $X=33470 $Y=405 $D=0
M23 4 3 VSS VSS N L=1.8e-07 W=9.4e-07 $X=35040 $Y=405 $D=0
M24 VDD 4 3 VDD P L=1.8e-07 W=1.095e-06 $X=620 $Y=2420 $D=16
M25 VDD 4 VDD VDD P L=9.9e-07 W=1.095e-06 $X=1340 $Y=2420 $D=16
M26 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=2870 $Y=2205 $D=16
M27 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=4400 $Y=2205 $D=16
M28 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=5930 $Y=2205 $D=16
M29 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=7460 $Y=2205 $D=16
M30 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=8990 $Y=2205 $D=16
M31 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=10520 $Y=2205 $D=16
M32 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=12050 $Y=2205 $D=16
M33 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=13580 $Y=2205 $D=16
M34 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=15110 $Y=2205 $D=16
M35 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=16640 $Y=2205 $D=16
M36 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=18170 $Y=2205 $D=16
M37 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=19700 $Y=2205 $D=16
M38 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=21230 $Y=2205 $D=16
M39 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=22760 $Y=2205 $D=16
M40 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=24290 $Y=2205 $D=16
M41 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=25820 $Y=2205 $D=16
M42 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=27350 $Y=2205 $D=16
M43 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=28880 $Y=2205 $D=16
M44 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=30410 $Y=2205 $D=16
M45 VDD 4 VDD VDD P L=9.9e-07 W=1.31e-06 $X=31940 $Y=2205 $D=16
M46 VDD 4 VDD VDD P L=9.9e-07 W=1.095e-06 $X=33470 $Y=2420 $D=16
M47 3 4 VDD VDD P L=1.8e-07 W=1.095e-06 $X=35040 $Y=2420 $D=16
.ENDS
***************************************
.SUBCKT ICV_46 1 2
** N=2 EP=2 IP=4 FDC=54
*.SEEDPROM
X0 1 2 DCAP8BWP7T $T=35840 0 0 0 $X=35550 $Y=-235
X1 2 1 DCAP64BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_36
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_47 1 2
** N=2 EP=2 IP=4 FDC=54
*.SEEDPROM
X0 1 2 ICV_46 $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT DCAP32BWP7T VDD VSS
** N=4 EP=2 IP=0 FDC=24
*.SEEDPROM
M0 VSS 3 4 VSS N L=1.8e-07 W=9.4e-07 $X=620 $Y=405 $D=0
M1 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=1340 $Y=405 $D=0
M2 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=2915 $Y=405 $D=0
M3 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=4490 $Y=405 $D=0
M4 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=6065 $Y=405 $D=0
M5 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=7640 $Y=405 $D=0
M6 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=9215 $Y=405 $D=0
M7 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=10790 $Y=405 $D=0
M8 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=12365 $Y=405 $D=0
M9 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=13940 $Y=405 $D=0
M10 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=15515 $Y=405 $D=0
M11 4 3 VSS VSS N L=1.8e-07 W=9.4e-07 $X=17120 $Y=405 $D=0
M12 VDD 4 3 VDD P L=1.8e-07 W=1.095e-06 $X=620 $Y=2420 $D=16
M13 VDD 4 VDD VDD P L=1.035e-06 W=1.095e-06 $X=1340 $Y=2420 $D=16
M14 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=2915 $Y=2205 $D=16
M15 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=4490 $Y=2205 $D=16
M16 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=6065 $Y=2205 $D=16
M17 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=7640 $Y=2205 $D=16
M18 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=9215 $Y=2205 $D=16
M19 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=10790 $Y=2205 $D=16
M20 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=12365 $Y=2205 $D=16
M21 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=13940 $Y=2205 $D=16
M22 VDD 4 VDD VDD P L=1.035e-06 W=1.095e-06 $X=15515 $Y=2420 $D=16
M23 3 4 VDD VDD P L=1.8e-07 W=1.095e-06 $X=17120 $Y=2420 $D=16
.ENDS
***************************************
.SUBCKT FA1D0BWP7T A B CI S VDD VSS CO
** N=18 EP=7 IP=0 FDC=28
*.SEEDPROM
M0 VSS A 8 VSS N L=1.8e-07 W=8.8e-07 $X=620 $Y=450 $D=0
M1 15 8 VSS VSS N L=1.8e-07 W=8.8e-07 $X=1340 $Y=450 $D=0
M2 9 11 15 VSS N L=1.8e-07 W=8.8e-07 $X=1940 $Y=450 $D=0
M3 8 B 9 VSS N L=1.8e-07 W=5e-07 $X=2700 $Y=830 $D=0
M4 VSS B 11 VSS N L=1.8e-07 W=4.25e-07 $X=4120 $Y=920 $D=0
M5 10 9 VSS VSS N L=1.8e-07 W=9.05e-07 $X=5040 $Y=440 $D=0
M6 14 10 11 VSS N L=1.8e-07 W=5.45e-07 $X=6460 $Y=780 $D=0
M7 12 9 14 VSS N L=1.8e-07 W=7e-07 $X=7180 $Y=555 $D=0
M8 13 10 12 VSS N L=1.8e-07 W=4.65e-07 $X=7900 $Y=790 $D=0
M9 16 9 13 VSS N L=1.8e-07 W=8.4e-07 $X=8620 $Y=415 $D=0
M10 VSS 12 16 VSS N L=1.8e-07 W=8.4e-07 $X=9140 $Y=415 $D=0
M11 12 CI VSS VSS N L=1.8e-07 W=8.4e-07 $X=9940 $Y=415 $D=0
M12 VSS 13 S VSS N L=1.8e-07 W=5e-07 $X=11360 $Y=350 $D=0
M13 CO 14 VSS VSS N L=1.8e-07 W=5e-07 $X=12080 $Y=350 $D=0
M14 VDD A 8 VDD P L=1.8e-07 W=1.18e-06 $X=620 $Y=2250 $D=16
M15 17 8 VDD VDD P L=1.8e-07 W=1.18e-06 $X=1340 $Y=2250 $D=16
M16 9 B 17 VDD P L=1.8e-07 W=1.02e-06 $X=1940 $Y=2410 $D=16
M17 8 11 9 VDD P L=1.8e-07 W=7.25e-07 $X=2660 $Y=2415 $D=16
M18 VDD B 11 VDD P L=1.8e-07 W=6.55e-07 $X=4080 $Y=2730 $D=16
M19 10 9 VDD VDD P L=1.8e-07 W=1.275e-06 $X=4880 $Y=2215 $D=16
M20 14 9 11 VDD P L=1.8e-07 W=1.01e-06 $X=6270 $Y=2450 $D=16
M21 12 10 14 VDD P L=1.8e-07 W=1.035e-06 $X=6990 $Y=2235 $D=16
M22 13 9 12 VDD P L=1.8e-07 W=8.8e-07 $X=7710 $Y=2235 $D=16
M23 18 10 13 VDD P L=1.8e-07 W=1e-06 $X=8430 $Y=2235 $D=16
M24 VDD 12 18 VDD P L=1.8e-07 W=1.16e-06 $X=9030 $Y=2235 $D=16
M25 12 CI VDD VDD P L=1.8e-07 W=1e-06 $X=9665 $Y=2210 $D=16
M26 VDD 13 S VDD P L=1.8e-07 W=6.85e-07 $X=11360 $Y=2315 $D=16
M27 CO 14 VDD VDD P L=1.8e-07 W=6.85e-07 $X=12080 $Y=2315 $D=16
.ENDS
***************************************
.SUBCKT INVD1BWP7T I VSS VDD ZN
** N=4 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=840 $Y=345 $D=0
M1 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=840 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKBD0BWP7T I VSS VDD Z
** N=5 EP=4 IP=0 FDC=4
*.SEEDPROM
M0 VSS I 5 VSS N L=1.8e-07 W=4.2e-07 $X=620 $Y=445 $D=0
M1 Z 5 VSS VSS N L=1.8e-07 W=4.2e-07 $X=1440 $Y=445 $D=0
M2 VDD I 5 VDD P L=1.8e-07 W=1.27e-06 $X=620 $Y=2290 $D=16
M3 Z 5 VDD VDD P L=1.8e-07 W=1.13e-06 $X=1440 $Y=2430 $D=16
.ENDS
***************************************
.SUBCKT FILL2BWP7T
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT FILL64BWP7T
** N=67 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT FILL32BWP7T
** N=35 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ND2D1BWP7T A2 VSS ZN A1 VDD
** N=6 EP=5 IP=0 FDC=4
*.SEEDPROM
M0 6 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=660 $Y=345 $D=0
M1 ZN A1 6 VSS N L=1.8e-07 W=1e-06 $X=1300 $Y=345 $D=0
M2 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M3 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1380 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_44
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT INVD0BWP7T I VSS VDD ZN
** N=4 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 ZN I VSS VSS N L=1.8e-07 W=5e-07 $X=840 $Y=560 $D=0
M1 ZN I VDD VDD P L=1.8e-07 W=6.85e-07 $X=840 $Y=2575 $D=16
.ENDS
***************************************
.SUBCKT OAI21D0BWP7T A2 ZN A1 B VSS VDD
** N=8 EP=6 IP=0 FDC=6
*.SEEDPROM
M0 ZN A2 7 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=845 $D=0
M1 7 A1 ZN VSS N L=1.8e-07 W=5e-07 $X=1340 $Y=845 $D=0
M2 VSS B 7 VSS N L=1.8e-07 W=4.65e-07 $X=2060 $Y=880 $D=0
M3 8 A2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2770 $D=16
M4 ZN A1 8 VDD P L=1.8e-07 W=6.85e-07 $X=1250 $Y=2770 $D=16
M5 VDD B ZN VDD P L=1.8e-07 W=6.85e-07 $X=1975 $Y=2770 $D=16
.ENDS
***************************************
.SUBCKT FILL16BWP7T
** N=19 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ND3D0BWP7T A3 VSS A2 A1 VDD ZN
** N=8 EP=6 IP=0 FDC=6
*.SEEDPROM
M0 7 A3 VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=500 $D=0
M1 8 A2 7 VSS N L=1.8e-07 W=5e-07 $X=1245 $Y=500 $D=0
M2 ZN A1 8 VSS N L=1.8e-07 W=5e-07 $X=1870 $Y=500 $D=0
M3 ZN A3 VDD VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2735 $D=16
M4 VDD A2 ZN VDD P L=1.8e-07 W=6.85e-07 $X=1340 $Y=2735 $D=16
M5 ZN A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=2000 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT DCAP16BWP7T VSS VDD
** N=4 EP=2 IP=0 FDC=12
*.SEEDPROM
M0 VSS 4 VSS VSS N L=9.65e-07 W=9.4e-07 $X=620 $Y=405 $D=0
M1 VSS 4 VSS VSS N L=9.65e-07 W=9.4e-07 $X=2125 $Y=405 $D=0
M2 VSS 4 VSS VSS N L=9.65e-07 W=9.4e-07 $X=3630 $Y=405 $D=0
M3 VSS 4 VSS VSS N L=9.65e-07 W=9.4e-07 $X=5135 $Y=405 $D=0
M4 VSS 4 VSS VSS N L=9.65e-07 W=9.4e-07 $X=6640 $Y=405 $D=0
M5 3 4 VSS VSS N L=1.8e-07 W=9.4e-07 $X=8160 $Y=405 $D=0
M6 VDD 3 VDD VDD P L=9.65e-07 W=1.31e-06 $X=620 $Y=2205 $D=16
M7 VDD 3 VDD VDD P L=9.65e-07 W=1.31e-06 $X=2125 $Y=2205 $D=16
M8 VDD 3 VDD VDD P L=9.65e-07 W=1.31e-06 $X=3630 $Y=2205 $D=16
M9 VDD 3 VDD VDD P L=9.65e-07 W=1.31e-06 $X=5135 $Y=2205 $D=16
M10 VDD 3 VDD VDD P L=9.65e-07 W=1.095e-06 $X=6640 $Y=2420 $D=16
M11 4 3 VDD VDD P L=1.8e-07 W=1.095e-06 $X=8160 $Y=2420 $D=16
.ENDS
***************************************
.SUBCKT FILL4BWP7T
** N=7 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT NR3D1BWP7T A1 VSS A2 A3 ZN VDD
** N=10 EP=6 IP=0 FDC=9
*.SEEDPROM
M0 ZN A3 VSS VSS N L=1.8e-07 W=1e-06 $X=640 $Y=345 $D=0
M1 VSS A2 ZN VSS N L=1.8e-07 W=1e-06 $X=1360 $Y=345 $D=0
M2 ZN A1 VSS VSS N L=1.8e-07 W=1e-06 $X=2160 $Y=345 $D=0
M3 7 A3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=640 $Y=2205 $D=16
M4 8 A2 7 VDD P L=1.8e-07 W=1.37e-06 $X=1230 $Y=2205 $D=16
M5 ZN A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=1820 $Y=2205 $D=16
M6 9 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2540 $Y=2205 $D=16
M7 10 A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=3095 $Y=2205 $D=16
M8 VDD A3 10 VDD P L=1.8e-07 W=1.37e-06 $X=3650 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT MAOI222D1BWP7T A C VSS VDD B ZN
** N=10 EP=6 IP=0 FDC=10
*.SEEDPROM
M0 ZN A 8 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 9 A ZN VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 VSS B 9 VSS N L=1.8e-07 W=1e-06 $X=1940 $Y=345 $D=0
M3 8 C VSS VSS N L=1.8e-07 W=1e-06 $X=2960 $Y=345 $D=0
M4 ZN B 8 VSS N L=1.8e-07 W=1e-06 $X=3680 $Y=345 $D=0
M5 ZN A 7 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M6 10 A ZN VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M7 VDD B 10 VDD P L=1.8e-07 W=1.37e-06 $X=2070 $Y=2205 $D=16
M8 7 C VDD VDD P L=1.8e-07 W=1.37e-06 $X=2960 $Y=2205 $D=16
M9 ZN B 7 VDD P L=1.8e-07 W=1.37e-06 $X=3680 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AOI21D1BWP7T A1 A2 VSS B ZN VDD
** N=8 EP=6 IP=0 FDC=6
*.SEEDPROM
M0 8 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=760 $Y=345 $D=0
M1 VSS A2 8 VSS N L=1.8e-07 W=1e-06 $X=1480 $Y=345 $D=0
M2 ZN B VSS VSS N L=1.8e-07 W=1e-06 $X=2200 $Y=345 $D=0
M3 ZN A1 7 VDD P L=1.8e-07 W=1.37e-06 $X=760 $Y=2205 $D=16
M4 7 A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1480 $Y=2205 $D=16
M5 VDD B 7 VDD P L=1.8e-07 W=1.37e-06 $X=2200 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INVD2BWP7T I ZN VDD VSS
** N=4 EP=4 IP=0 FDC=4
*.SEEDPROM
M0 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=670 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=1390 $Y=345 $D=0
M2 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=670 $Y=2205 $D=16
M3 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1390 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT FILL8BWP7T
** N=11 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT DFQD0BWP7T CP D VSS VDD Q
** N=16 EP=5 IP=0 FDC=24
*.SEEDPROM
M0 VSS CP 6 VSS N L=1.8e-07 W=5e-07 $X=640 $Y=840 $D=0
M1 9 6 VSS VSS N L=1.8e-07 W=5e-07 $X=1240 $Y=840 $D=0
M2 13 6 VSS VSS N L=1.8e-07 W=9.4e-07 $X=2665 $Y=405 $D=0
M3 7 D 13 VSS N L=1.8e-07 W=9.4e-07 $X=3135 $Y=405 $D=0
M4 14 9 7 VSS N L=1.8e-07 W=4.2e-07 $X=3990 $Y=895 $D=0
M5 VSS 8 14 VSS N L=1.8e-07 W=4.2e-07 $X=4485 $Y=895 $D=0
M6 8 7 VSS VSS N L=1.8e-07 W=5.4e-07 $X=5285 $Y=775 $D=0
M7 11 9 8 VSS N L=1.8e-07 W=9.1e-07 $X=6005 $Y=405 $D=0
M8 10 6 11 VSS N L=1.8e-07 W=4.2e-07 $X=6725 $Y=895 $D=0
M9 VSS 12 10 VSS N L=1.8e-07 W=4.2e-07 $X=7445 $Y=895 $D=0
M10 12 11 VSS VSS N L=1.8e-07 W=5e-07 $X=8300 $Y=430 $D=0
M11 Q 12 VSS VSS N L=1.8e-07 W=5e-07 $X=9840 $Y=430 $D=0
M12 VDD CP 6 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2345 $D=16
M13 9 6 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1240 $Y=2345 $D=16
M14 15 9 VDD VDD P L=1.8e-07 W=9.2e-07 $X=2705 $Y=2205 $D=16
M15 7 D 15 VDD P L=1.8e-07 W=9.2e-07 $X=3205 $Y=2205 $D=16
M16 16 6 7 VDD P L=1.8e-07 W=4.2e-07 $X=3985 $Y=2705 $D=16
M17 VDD 8 16 VDD P L=1.8e-07 W=4.2e-07 $X=4485 $Y=2705 $D=16
M18 8 7 VDD VDD P L=1.8e-07 W=9.6e-07 $X=5285 $Y=2175 $D=16
M19 11 6 8 VDD P L=1.8e-07 W=1.34e-06 $X=6005 $Y=2175 $D=16
M20 10 9 11 VDD P L=1.8e-07 W=4.2e-07 $X=6725 $Y=2470 $D=16
M21 VDD 12 10 VDD P L=1.8e-07 W=4.2e-07 $X=7485 $Y=2205 $D=16
M22 12 11 VDD VDD P L=1.8e-07 W=6.85e-07 $X=8300 $Y=2890 $D=16
M23 Q 12 VDD VDD P L=1.8e-07 W=6.85e-07 $X=9840 $Y=2670 $D=16
.ENDS
***************************************
.SUBCKT INVD4BWP7T I ZN VSS VDD
** N=4 EP=4 IP=0 FDC=8
*.SEEDPROM
M0 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=765 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=1485 $Y=345 $D=0
M2 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=2275 $Y=345 $D=0
M3 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=2995 $Y=345 $D=0
M4 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=765 $Y=2205 $D=16
M5 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1485 $Y=2205 $D=16
M6 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=2275 $Y=2205 $D=16
M7 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=2995 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR3D0BWP7T A3 VSS VDD A2 A1 ZN
** N=8 EP=6 IP=0 FDC=6
*.SEEDPROM
M0 ZN A3 VSS VSS N L=1.8e-07 W=5e-07 $X=625 $Y=770 $D=0
M1 VSS A2 ZN VSS N L=1.8e-07 W=5e-07 $X=1345 $Y=770 $D=0
M2 ZN A1 VSS VSS N L=1.8e-07 W=5e-07 $X=2000 $Y=770 $D=0
M3 7 A3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=625 $Y=2205 $D=16
M4 8 A2 7 VDD P L=1.8e-07 W=1.37e-06 $X=1225 $Y=2205 $D=16
M5 ZN A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=1825 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AOI21D2BWP7T B VDD ZN A1 A2 VSS
** N=9 EP=6 IP=0 FDC=12
*.SEEDPROM
M0 ZN B VSS VSS N L=1.8e-07 W=1e-06 $X=625 $Y=345 $D=0
M1 VSS B ZN VSS N L=1.8e-07 W=1e-06 $X=1345 $Y=345 $D=0
M2 8 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=2145 $Y=345 $D=0
M3 ZN A1 8 VSS N L=1.8e-07 W=1e-06 $X=2800 $Y=345 $D=0
M4 9 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=3520 $Y=345 $D=0
M5 VSS A2 9 VSS N L=1.8e-07 W=1e-06 $X=4240 $Y=345 $D=0
M6 VDD B 7 VDD P L=1.8e-07 W=1.37e-06 $X=625 $Y=2205 $D=16
M7 7 B VDD VDD P L=1.8e-07 W=1.37e-06 $X=1345 $Y=2205 $D=16
M8 ZN A2 7 VDD P L=1.8e-07 W=1.37e-06 $X=2080 $Y=2205 $D=16
M9 7 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2800 $Y=2205 $D=16
M10 ZN A1 7 VDD P L=1.8e-07 W=1.37e-06 $X=3520 $Y=2205 $D=16
M11 7 A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4240 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AOI21D0BWP7T A2 ZN A1 B VSS VDD
** N=8 EP=6 IP=0 FDC=6
*.SEEDPROM
M0 8 A2 VSS VSS N L=1.8e-07 W=5e-07 $X=630 $Y=460 $D=0
M1 ZN A1 8 VSS N L=1.8e-07 W=5e-07 $X=1250 $Y=460 $D=0
M2 VSS B ZN VSS N L=1.8e-07 W=5e-07 $X=1975 $Y=460 $D=0
M3 ZN A2 7 VDD P L=1.8e-07 W=6.85e-07 $X=630 $Y=2275 $D=16
M4 7 A1 ZN VDD P L=1.8e-07 W=6.85e-07 $X=1355 $Y=2275 $D=16
M5 VDD B 7 VDD P L=1.8e-07 W=6.85e-07 $X=2075 $Y=2275 $D=16
.ENDS
***************************************
.SUBCKT BUFFD0BWP7T I VSS VDD Z
** N=5 EP=4 IP=0 FDC=4
*.SEEDPROM
M0 VSS I 5 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=555 $D=0
M1 Z 5 VSS VSS N L=1.8e-07 W=5e-07 $X=1420 $Y=555 $D=0
M2 VDD I 5 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2850 $D=16
M3 Z 5 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1420 $Y=2850 $D=16
.ENDS
***************************************
.SUBCKT AN2D1BWP7T A1 A2 VSS VDD Z
** N=7 EP=5 IP=0 FDC=6
*.SEEDPROM
M0 7 A1 6 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=345 $D=0
M1 VSS A2 7 VSS N L=1.8e-07 W=5e-07 $X=1205 $Y=345 $D=0
M2 Z 6 VSS VSS N L=1.8e-07 W=1e-06 $X=2000 $Y=345 $D=0
M3 6 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=520 $Y=2205 $D=16
M4 VDD A2 6 VDD P L=1.8e-07 W=6.85e-07 $X=1240 $Y=2205 $D=16
M5 Z 6 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2000 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_61 1 2
** N=2 EP=2 IP=4 FDC=16
*.SEEDPROM
X0 1 2 DCAP4BWP7T $T=8960 0 0 0 $X=8670 $Y=-235
X1 1 2 DCAP16BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT XOR3D0BWP7T A2 A1 A3 VDD VSS Z
** N=16 EP=6 IP=0 FDC=22
*.SEEDPROM
M0 VSS A2 7 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=480 $D=0
M1 13 8 VSS VSS N L=1.8e-07 W=5e-07 $X=1405 $Y=845 $D=0
M2 9 A2 13 VSS N L=1.8e-07 W=5e-07 $X=2025 $Y=480 $D=0
M3 8 7 9 VSS N L=1.8e-07 W=5e-07 $X=2825 $Y=480 $D=0
M4 VSS A1 8 VSS N L=1.8e-07 W=5e-07 $X=3585 $Y=480 $D=0
M5 VSS 9 10 VSS N L=1.8e-07 W=5e-07 $X=5115 $Y=460 $D=0
M6 14 11 VSS VSS N L=1.8e-07 W=5e-07 $X=5915 $Y=845 $D=0
M7 12 10 14 VSS N L=1.8e-07 W=5e-07 $X=6345 $Y=845 $D=0
M8 11 9 12 VSS N L=1.8e-07 W=5e-07 $X=7205 $Y=440 $D=0
M9 VSS A3 11 VSS N L=1.8e-07 W=5e-07 $X=7965 $Y=440 $D=0
M10 Z 12 VSS VSS N L=1.8e-07 W=5e-07 $X=8715 $Y=440 $D=0
M11 VDD A2 7 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2795 $D=16
M12 15 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1405 $Y=2425 $D=16
M13 9 7 15 VDD P L=1.8e-07 W=6.85e-07 $X=1985 $Y=2425 $D=16
M14 8 A2 9 VDD P L=1.8e-07 W=6.85e-07 $X=2785 $Y=2425 $D=16
M15 VDD A1 8 VDD P L=1.8e-07 W=6.85e-07 $X=3545 $Y=2425 $D=16
M16 VDD 9 10 VDD P L=1.8e-07 W=6.85e-07 $X=5115 $Y=2815 $D=16
M17 16 11 VDD VDD P L=1.8e-07 W=6.85e-07 $X=5915 $Y=2445 $D=16
M18 12 9 16 VDD P L=1.8e-07 W=6.85e-07 $X=6425 $Y=2445 $D=16
M19 11 10 12 VDD P L=1.8e-07 W=6.85e-07 $X=7165 $Y=2205 $D=16
M20 VDD A3 11 VDD P L=1.8e-07 W=6.85e-07 $X=7915 $Y=2205 $D=16
M21 Z 12 VDD VDD P L=1.8e-07 W=6.85e-07 $X=8715 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT XNR3D0BWP7T A2 A1 A3 VDD VSS ZN
** N=16 EP=6 IP=0 FDC=22
*.SEEDPROM
M0 VSS A2 7 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=845 $D=0
M1 13 8 VSS VSS N L=1.8e-07 W=5e-07 $X=1500 $Y=845 $D=0
M2 9 7 13 VSS N L=1.8e-07 W=5e-07 $X=2045 $Y=845 $D=0
M3 8 A2 9 VSS N L=1.8e-07 W=5e-07 $X=2825 $Y=845 $D=0
M4 VSS A1 8 VSS N L=1.8e-07 W=7.05e-07 $X=3545 $Y=640 $D=0
M5 VSS 9 10 VSS N L=1.8e-07 W=5e-07 $X=5115 $Y=460 $D=0
M6 14 11 VSS VSS N L=1.8e-07 W=5e-07 $X=5915 $Y=845 $D=0
M7 12 10 14 VSS N L=1.8e-07 W=5e-07 $X=6345 $Y=845 $D=0
M8 11 9 12 VSS N L=1.8e-07 W=5e-07 $X=7205 $Y=440 $D=0
M9 VSS A3 11 VSS N L=1.8e-07 W=5e-07 $X=7965 $Y=440 $D=0
M10 ZN 12 VSS VSS N L=1.8e-07 W=5e-07 $X=8720 $Y=440 $D=0
M11 VDD A2 7 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2645 $D=16
M12 15 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1420 $Y=2435 $D=16
M13 9 A2 15 VDD P L=1.8e-07 W=6.85e-07 $X=1900 $Y=2435 $D=16
M14 8 7 9 VDD P L=1.8e-07 W=6.85e-07 $X=2745 $Y=2435 $D=16
M15 VDD A1 8 VDD P L=1.8e-07 W=6.85e-07 $X=3545 $Y=2435 $D=16
M16 VDD 9 10 VDD P L=1.8e-07 W=6.85e-07 $X=5115 $Y=2815 $D=16
M17 16 11 VDD VDD P L=1.8e-07 W=6.85e-07 $X=5915 $Y=2445 $D=16
M18 12 9 16 VDD P L=1.8e-07 W=6.85e-07 $X=6425 $Y=2445 $D=16
M19 11 10 12 VDD P L=1.8e-07 W=6.85e-07 $X=7145 $Y=2445 $D=16
M20 VDD A3 11 VDD P L=1.8e-07 W=6.85e-07 $X=7905 $Y=2205 $D=16
M21 ZN 12 VDD VDD P L=1.8e-07 W=6.85e-07 $X=8720 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OAI22D1BWP7T B1 B2 VSS A2 VDD ZN A1
** N=10 EP=7 IP=0 FDC=8
*.SEEDPROM
M0 VSS B1 8 VSS N L=1.8e-07 W=1e-06 $X=640 $Y=345 $D=0
M1 8 B2 VSS VSS N L=1.8e-07 W=1e-06 $X=1440 $Y=345 $D=0
M2 ZN A2 8 VSS N L=1.8e-07 W=1e-06 $X=2180 $Y=345 $D=0
M3 8 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=3120 $Y=345 $D=0
M4 9 B1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=640 $Y=2205 $D=16
M5 VDD B2 9 VDD P L=1.8e-07 W=1.37e-06 $X=1440 $Y=2205 $D=16
M6 10 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2420 $Y=2205 $D=16
M7 ZN A1 10 VDD P L=1.8e-07 W=1.37e-06 $X=3120 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IOA21D0BWP7T A1 A2 VSS ZN B VDD
** N=9 EP=6 IP=0 FDC=8
*.SEEDPROM
M0 8 A1 7 VSS N L=1.8e-07 W=4.2e-07 $X=625 $Y=440 $D=0
M1 VSS A2 8 VSS N L=1.8e-07 W=4.2e-07 $X=1205 $Y=440 $D=0
M2 9 7 VSS VSS N L=1.8e-07 W=5e-07 $X=1945 $Y=360 $D=0
M3 ZN B 9 VSS N L=1.8e-07 W=5e-07 $X=2560 $Y=360 $D=0
M4 7 A1 VDD VDD P L=1.8e-07 W=4.2e-07 $X=465 $Y=2500 $D=16
M5 VDD A2 7 VDD P L=1.8e-07 W=4.2e-07 $X=1185 $Y=2500 $D=16
M6 ZN 7 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1840 $Y=2500 $D=16
M7 VDD B ZN VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2500 $D=16
.ENDS
***************************************
.SUBCKT OAI211D0BWP7T C VSS B A1 VDD A2 ZN
** N=10 EP=7 IP=0 FDC=8
*.SEEDPROM
M0 8 C VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=680 $D=0
M1 9 B 8 VSS N L=1.8e-07 W=5e-07 $X=1115 $Y=680 $D=0
M2 ZN A1 9 VSS N L=1.8e-07 W=5e-07 $X=1820 $Y=680 $D=0
M3 9 A2 ZN VSS N L=1.8e-07 W=5e-07 $X=2560 $Y=680 $D=0
M4 ZN C VDD VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2830 $D=16
M5 VDD B ZN VDD P L=1.8e-07 W=6.85e-07 $X=1340 $Y=2830 $D=16
M6 10 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=2060 $Y=2830 $D=16
M7 ZN A2 10 VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2830 $D=16
.ENDS
***************************************
.SUBCKT AO22D0BWP7T B2 A1 A2 B1 VSS VDD Z
** N=11 EP=7 IP=0 FDC=10
*.SEEDPROM
M0 10 B2 VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=460 $D=0
M1 8 B1 10 VSS N L=1.8e-07 W=5e-07 $X=1115 $Y=460 $D=0
M2 11 A1 8 VSS N L=1.8e-07 W=5e-07 $X=1915 $Y=460 $D=0
M3 VSS A2 11 VSS N L=1.8e-07 W=5e-07 $X=2475 $Y=460 $D=0
M4 Z 8 VSS VSS N L=1.8e-07 W=5e-07 $X=3675 $Y=460 $D=0
M5 9 B2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2670 $D=16
M6 8 A1 9 VDD P L=1.8e-07 W=6.85e-07 $X=1415 $Y=2670 $D=16
M7 9 A2 8 VDD P L=1.8e-07 W=6.85e-07 $X=2235 $Y=2670 $D=16
M8 VDD B1 9 VDD P L=1.8e-07 W=6.85e-07 $X=2955 $Y=2670 $D=16
M9 Z 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=3675 $Y=2670 $D=16
.ENDS
***************************************
.SUBCKT MAOI222D2BWP7T A C B ZN VSS VDD
** N=12 EP=6 IP=0 FDC=16
*.SEEDPROM
M0 9 A 8 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 11 A 9 VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 VSS B 11 VSS N L=1.8e-07 W=1e-06 $X=1940 $Y=345 $D=0
M3 8 C VSS VSS N L=1.8e-07 W=1e-06 $X=2740 $Y=345 $D=0
M4 9 B 8 VSS N L=1.8e-07 W=1e-06 $X=3460 $Y=345 $D=0
M5 VSS 9 10 VSS N L=1.8e-07 W=1e-06 $X=5015 $Y=345 $D=0
M6 ZN 10 VSS VSS N L=1.8e-07 W=1e-06 $X=5735 $Y=345 $D=0
M7 VSS 10 ZN VSS N L=1.8e-07 W=1e-06 $X=6455 $Y=345 $D=0
M8 9 A 7 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M9 12 A 9 VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M10 VDD B 12 VDD P L=1.8e-07 W=1.37e-06 $X=1940 $Y=2205 $D=16
M11 7 C VDD VDD P L=1.8e-07 W=1.37e-06 $X=2740 $Y=2205 $D=16
M12 9 B 7 VDD P L=1.8e-07 W=1.37e-06 $X=3460 $Y=2205 $D=16
M13 VDD 9 10 VDD P L=1.8e-07 W=1.37e-06 $X=5015 $Y=2205 $D=16
M14 ZN 10 VDD VDD P L=1.8e-07 W=1.37e-06 $X=5735 $Y=2205 $D=16
M15 VDD 10 ZN VDD P L=1.8e-07 W=1.37e-06 $X=6455 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT DFQD1BWP7T CP D VSS VDD Q
** N=16 EP=5 IP=0 FDC=24
*.SEEDPROM
M0 VSS CP 6 VSS N L=1.8e-07 W=5e-07 $X=640 $Y=840 $D=0
M1 9 6 VSS VSS N L=1.8e-07 W=5e-07 $X=1240 $Y=840 $D=0
M2 13 6 VSS VSS N L=1.8e-07 W=9.4e-07 $X=2665 $Y=405 $D=0
M3 7 D 13 VSS N L=1.8e-07 W=9.4e-07 $X=3135 $Y=405 $D=0
M4 14 9 7 VSS N L=1.8e-07 W=4.2e-07 $X=3990 $Y=895 $D=0
M5 VSS 8 14 VSS N L=1.8e-07 W=4.2e-07 $X=4485 $Y=895 $D=0
M6 8 7 VSS VSS N L=1.8e-07 W=5.4e-07 $X=5285 $Y=775 $D=0
M7 11 9 8 VSS N L=1.8e-07 W=9.1e-07 $X=6005 $Y=405 $D=0
M8 10 6 11 VSS N L=1.8e-07 W=4.2e-07 $X=6725 $Y=895 $D=0
M9 VSS 12 10 VSS N L=1.8e-07 W=4.2e-07 $X=7445 $Y=895 $D=0
M10 12 11 VSS VSS N L=1.8e-07 W=1e-06 $X=8300 $Y=345 $D=0
M11 Q 12 VSS VSS N L=1.8e-07 W=1e-06 $X=9840 $Y=345 $D=0
M12 VDD CP 6 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2345 $D=16
M13 9 6 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1240 $Y=2345 $D=16
M14 15 9 VDD VDD P L=1.8e-07 W=9.2e-07 $X=2705 $Y=2205 $D=16
M15 7 D 15 VDD P L=1.8e-07 W=9.2e-07 $X=3205 $Y=2205 $D=16
M16 16 6 7 VDD P L=1.8e-07 W=4.2e-07 $X=3985 $Y=2705 $D=16
M17 VDD 8 16 VDD P L=1.8e-07 W=4.2e-07 $X=4485 $Y=2705 $D=16
M18 8 7 VDD VDD P L=1.8e-07 W=9.6e-07 $X=5285 $Y=2175 $D=16
M19 11 6 8 VDD P L=1.8e-07 W=1.34e-06 $X=6005 $Y=2175 $D=16
M20 10 9 11 VDD P L=1.8e-07 W=4.2e-07 $X=6725 $Y=2470 $D=16
M21 VDD 12 10 VDD P L=1.8e-07 W=4.2e-07 $X=7485 $Y=2205 $D=16
M22 12 11 VDD VDD P L=1.8e-07 W=1.37e-06 $X=8300 $Y=2205 $D=16
M23 Q 12 VDD VDD P L=1.8e-07 W=1.37e-06 $X=9840 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT MOAI22D0BWP7T B1 B2 VSS VDD A1 ZN A2
** N=11 EP=7 IP=0 FDC=10
*.SEEDPROM
M0 9 B1 8 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=610 $D=0
M1 VSS B2 9 VSS N L=1.8e-07 W=5e-07 $X=1050 $Y=610 $D=0
M2 10 8 VSS VSS N L=1.8e-07 W=5e-07 $X=1850 $Y=610 $D=0
M3 ZN A1 10 VSS N L=1.8e-07 W=5e-07 $X=2560 $Y=845 $D=0
M4 10 A2 ZN VSS N L=1.8e-07 W=5e-07 $X=3280 $Y=845 $D=0
M5 8 B1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=460 $Y=2390 $D=16
M6 VDD B2 8 VDD P L=1.8e-07 W=6.85e-07 $X=1180 $Y=2390 $D=16
M7 ZN 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1980 $Y=2390 $D=16
M8 11 A1 ZN VDD P L=1.8e-07 W=6.85e-07 $X=2700 $Y=2390 $D=16
M9 VDD A2 11 VDD P L=1.8e-07 W=6.85e-07 $X=3280 $Y=2390 $D=16
.ENDS
***************************************
.SUBCKT XNR4D0BWP7T A4 A3 ZN A2 A1 VSS VDD
** N=21 EP=7 IP=0 FDC=30
*.SEEDPROM
M0 VSS A4 8 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=500 $D=0
M1 16 9 VSS VSS N L=1.8e-07 W=5e-07 $X=1445 $Y=835 $D=0
M2 10 A4 16 VSS N L=1.8e-07 W=5e-07 $X=1925 $Y=835 $D=0
M3 9 8 10 VSS N L=1.8e-07 W=5e-07 $X=2645 $Y=835 $D=0
M4 VSS A3 9 VSS N L=1.8e-07 W=5e-07 $X=3425 $Y=835 $D=0
M5 VSS 10 11 VSS N L=1.8e-07 W=5e-07 $X=4980 $Y=775 $D=0
M6 17 13 VSS VSS N L=1.8e-07 W=5e-07 $X=5700 $Y=775 $D=0
M7 12 10 17 VSS N L=1.8e-07 W=5e-07 $X=6180 $Y=775 $D=0
M8 13 11 12 VSS N L=1.8e-07 W=5e-07 $X=6900 $Y=775 $D=0
M9 VSS 12 ZN VSS N L=1.8e-07 W=5e-07 $X=8320 $Y=630 $D=0
M10 14 A2 VSS VSS N L=1.8e-07 W=5e-07 $X=9120 $Y=630 $D=0
M11 13 15 14 VSS N L=1.8e-07 W=5e-07 $X=9885 $Y=775 $D=0
M12 18 A1 13 VSS N L=1.8e-07 W=5e-07 $X=10605 $Y=775 $D=0
M13 VSS 14 18 VSS N L=1.8e-07 W=5e-07 $X=11320 $Y=775 $D=0
M14 15 A1 VSS VSS N L=1.8e-07 W=5e-07 $X=12080 $Y=595 $D=0
M15 VDD A4 8 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2710 $D=16
M16 19 9 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1380 $Y=2460 $D=16
M17 10 8 19 VDD P L=1.8e-07 W=6.85e-07 $X=1925 $Y=2460 $D=16
M18 9 A4 10 VDD P L=1.8e-07 W=6.85e-07 $X=2645 $Y=2460 $D=16
M19 VDD A3 9 VDD P L=1.8e-07 W=6.85e-07 $X=3425 $Y=2205 $D=16
M20 VDD 10 11 VDD P L=1.8e-07 W=6.85e-07 $X=4980 $Y=2370 $D=16
M21 20 13 VDD VDD P L=1.8e-07 W=6.85e-07 $X=5700 $Y=2370 $D=16
M22 12 11 20 VDD P L=1.8e-07 W=6.85e-07 $X=6180 $Y=2370 $D=16
M23 13 10 12 VDD P L=1.8e-07 W=6.85e-07 $X=6900 $Y=2370 $D=16
M24 VDD 12 ZN VDD P L=1.8e-07 W=6.85e-07 $X=8320 $Y=2205 $D=16
M25 14 A2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=9120 $Y=2205 $D=16
M26 13 A1 14 VDD P L=1.8e-07 W=6.85e-07 $X=9885 $Y=2385 $D=16
M27 21 15 13 VDD P L=1.8e-07 W=6.85e-07 $X=10605 $Y=2385 $D=16
M28 VDD 14 21 VDD P L=1.8e-07 W=6.85e-07 $X=11290 $Y=2385 $D=16
M29 15 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=12080 $Y=2720 $D=16
.ENDS
***************************************
.SUBCKT BUFFD12BWP7T I Z VSS VDD
** N=5 EP=4 IP=0 FDC=32
*.SEEDPROM
M0 5 I VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 5 I VSS VSS N L=1.8e-07 W=1e-06 $X=2060 $Y=345 $D=0
M3 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=2780 $Y=345 $D=0
M4 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=3500 $Y=345 $D=0
M5 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=4220 $Y=345 $D=0
M6 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=4940 $Y=345 $D=0
M7 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=5660 $Y=345 $D=0
M8 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=6400 $Y=345 $D=0
M9 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=7120 $Y=345 $D=0
M10 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=7850 $Y=345 $D=0
M11 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=8570 $Y=345 $D=0
M12 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=9300 $Y=345 $D=0
M13 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=10020 $Y=345 $D=0
M14 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=10740 $Y=345 $D=0
M15 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=11500 $Y=345 $D=0
M16 5 I VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M17 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M18 5 I VDD VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M19 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M20 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3500 $Y=2205 $D=16
M21 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=4220 $Y=2205 $D=16
M22 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4940 $Y=2205 $D=16
M23 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=5660 $Y=2205 $D=16
M24 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=6400 $Y=2205 $D=16
M25 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=7120 $Y=2205 $D=16
M26 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=7850 $Y=2205 $D=16
M27 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=8570 $Y=2205 $D=16
M28 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=9300 $Y=2205 $D=16
M29 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=10020 $Y=2205 $D=16
M30 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=10740 $Y=2205 $D=16
M31 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=11500 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OAI22D2BWP7T B1 VSS B2 ZN A1 A2 VDD
** N=12 EP=7 IP=0 FDC=16
*.SEEDPROM
M0 VSS B2 8 VSS N L=1.8e-07 W=1e-06 $X=630 $Y=345 $D=0
M1 8 B1 VSS VSS N L=1.8e-07 W=1e-06 $X=1400 $Y=345 $D=0
M2 VSS B1 8 VSS N L=1.8e-07 W=1e-06 $X=2120 $Y=345 $D=0
M3 8 B2 VSS VSS N L=1.8e-07 W=1e-06 $X=2920 $Y=345 $D=0
M4 ZN A2 8 VSS N L=1.8e-07 W=1e-06 $X=3680 $Y=345 $D=0
M5 8 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=4420 $Y=345 $D=0
M6 ZN A1 8 VSS N L=1.8e-07 W=1e-06 $X=5140 $Y=345 $D=0
M7 8 A2 ZN VSS N L=1.8e-07 W=1e-06 $X=5860 $Y=345 $D=0
M8 9 B2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=630 $Y=2205 $D=16
M9 ZN B1 9 VDD P L=1.8e-07 W=1.37e-06 $X=1400 $Y=2205 $D=16
M10 10 B1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2120 $Y=2205 $D=16
M11 VDD B2 10 VDD P L=1.8e-07 W=1.37e-06 $X=2760 $Y=2205 $D=16
M12 11 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3720 $Y=2205 $D=16
M13 ZN A1 11 VDD P L=1.8e-07 W=1.37e-06 $X=4320 $Y=2205 $D=16
M14 12 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=5080 $Y=2205 $D=16
M15 VDD A2 12 VDD P L=1.8e-07 W=1.37e-06 $X=5680 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT XOR4D0BWP7T A4 A3 Z A2 A1 VSS VDD
** N=21 EP=7 IP=0 FDC=30
*.SEEDPROM
M0 VSS A4 8 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=600 $D=0
M1 16 9 VSS VSS N L=1.8e-07 W=5e-07 $X=1380 $Y=775 $D=0
M2 10 A4 16 VSS N L=1.8e-07 W=5e-07 $X=2010 $Y=775 $D=0
M3 9 8 10 VSS N L=1.8e-07 W=5e-07 $X=2730 $Y=775 $D=0
M4 VSS A3 9 VSS N L=1.8e-07 W=5e-07 $X=3510 $Y=585 $D=0
M5 VSS 10 11 VSS N L=1.8e-07 W=5e-07 $X=4930 $Y=845 $D=0
M6 17 13 VSS VSS N L=1.8e-07 W=5e-07 $X=5650 $Y=845 $D=0
M7 12 11 17 VSS N L=1.8e-07 W=5e-07 $X=6130 $Y=845 $D=0
M8 13 10 12 VSS N L=1.8e-07 W=5e-07 $X=6890 $Y=440 $D=0
M9 VSS 12 Z VSS N L=1.8e-07 W=5e-07 $X=8320 $Y=630 $D=0
M10 14 A2 VSS VSS N L=1.8e-07 W=5e-07 $X=9120 $Y=630 $D=0
M11 13 15 14 VSS N L=1.8e-07 W=5e-07 $X=9885 $Y=775 $D=0
M12 18 A1 13 VSS N L=1.8e-07 W=5e-07 $X=10605 $Y=775 $D=0
M13 VSS 14 18 VSS N L=1.8e-07 W=5e-07 $X=11320 $Y=775 $D=0
M14 15 A1 VSS VSS N L=1.8e-07 W=5e-07 $X=12080 $Y=595 $D=0
M15 VDD A4 8 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2675 $D=16
M16 19 9 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1380 $Y=2430 $D=16
M17 10 8 19 VDD P L=1.8e-07 W=6.85e-07 $X=2010 $Y=2430 $D=16
M18 9 A4 10 VDD P L=1.8e-07 W=6.85e-07 $X=2750 $Y=2430 $D=16
M19 VDD A3 9 VDD P L=1.8e-07 W=6.85e-07 $X=3470 $Y=2430 $D=16
M20 VDD 10 11 VDD P L=1.8e-07 W=6.85e-07 $X=4930 $Y=2405 $D=16
M21 20 13 VDD VDD P L=1.8e-07 W=6.85e-07 $X=5650 $Y=2405 $D=16
M22 12 10 20 VDD P L=1.8e-07 W=6.85e-07 $X=6140 $Y=2405 $D=16
M23 13 11 12 VDD P L=1.8e-07 W=6.85e-07 $X=6880 $Y=2405 $D=16
M24 VDD 12 Z VDD P L=1.8e-07 W=6.85e-07 $X=8320 $Y=2205 $D=16
M25 14 A2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=9120 $Y=2205 $D=16
M26 13 A1 14 VDD P L=1.8e-07 W=6.85e-07 $X=9885 $Y=2385 $D=16
M27 21 15 13 VDD P L=1.8e-07 W=6.85e-07 $X=10605 $Y=2385 $D=16
M28 VDD 14 21 VDD P L=1.8e-07 W=6.85e-07 $X=11290 $Y=2385 $D=16
M29 15 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=12080 $Y=2720 $D=16
.ENDS
***************************************
.SUBCKT CKND1BWP7T I VSS VDD ZN
** N=4 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 ZN I VSS VSS N L=1.8e-07 W=5.25e-07 $X=830 $Y=440 $D=0
M1 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=830 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IAO22D2BWP7T A2 A1 ZN B1 VSS B2 VDD
** N=12 EP=7 IP=0 FDC=14
*.SEEDPROM
M0 8 10 9 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS A2 8 VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 8 A1 VSS VSS N L=1.8e-07 W=1e-06 $X=2140 $Y=345 $D=0
M3 ZN 9 VSS VSS N L=1.8e-07 W=1e-06 $X=3490 $Y=345 $D=0
M4 VSS 9 ZN VSS N L=1.8e-07 W=1e-06 $X=4210 $Y=345 $D=0
M5 11 B1 VSS VSS N L=1.8e-07 W=5e-07 $X=4930 $Y=345 $D=0
M6 10 B2 11 VSS N L=1.8e-07 W=5e-07 $X=5360 $Y=345 $D=0
M7 9 10 VDD VDD P L=1.8e-07 W=1.37e-06 $X=685 $Y=2205 $D=16
M8 12 A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=1405 $Y=2205 $D=16
M9 VDD A1 12 VDD P L=1.8e-07 W=1.37e-06 $X=1965 $Y=2205 $D=16
M10 ZN 9 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2795 $Y=2205 $D=16
M11 VDD 9 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3840 $Y=2205 $D=16
M12 10 B1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=4640 $Y=2820 $D=16
M13 VDD B2 10 VDD P L=1.8e-07 W=6.85e-07 $X=5360 $Y=2820 $D=16
.ENDS
***************************************
.SUBCKT BUFFD1P5BWP7T I Z VSS VDD
** N=5 EP=4 IP=0 FDC=6
*.SEEDPROM
M0 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 VSS 5 Z VSS N L=1.8e-07 W=4.65e-07 $X=2060 $Y=880 $D=0
M3 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M4 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M5 VDD 5 Z VDD P L=1.8e-07 W=6.85e-07 $X=2060 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKND2BWP7T I ZN VDD VSS
** N=4 EP=4 IP=0 FDC=4
*.SEEDPROM
M0 ZN I VSS VSS N L=1.8e-07 W=5.25e-07 $X=670 $Y=440 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=5.25e-07 $X=1390 $Y=440 $D=0
M2 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=670 $Y=2205 $D=16
M3 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1390 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR2D0BWP7T A2 VDD A1 ZN VSS
** N=6 EP=5 IP=0 FDC=4
*.SEEDPROM
M0 ZN A2 VSS VSS N L=1.8e-07 W=5e-07 $X=660 $Y=500 $D=0
M1 VSS A1 ZN VSS N L=1.8e-07 W=5e-07 $X=1380 $Y=500 $D=0
M2 6 A2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=660 $Y=2735 $D=16
M3 ZN A1 6 VDD P L=1.8e-07 W=6.85e-07 $X=1260 $Y=2735 $D=16
.ENDS
***************************************
.SUBCKT AOI22D1BWP7T B1 B2 VDD A2 VSS A1 ZN
** N=10 EP=7 IP=0 FDC=8
*.SEEDPROM
M0 9 B1 ZN VSS N L=1.8e-07 W=1e-06 $X=640 $Y=345 $D=0
M1 VSS B2 9 VSS N L=1.8e-07 W=1e-06 $X=1440 $Y=345 $D=0
M2 10 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=2420 $Y=345 $D=0
M3 ZN A1 10 VSS N L=1.8e-07 W=1e-06 $X=3120 $Y=345 $D=0
M4 VDD B1 8 VDD P L=1.8e-07 W=1.37e-06 $X=640 $Y=2205 $D=16
M5 8 B2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1440 $Y=2205 $D=16
M6 ZN A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=2180 $Y=2205 $D=16
M7 8 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3120 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INVD3BWP7T I VSS VDD ZN
** N=4 EP=4 IP=0 FDC=6
*.SEEDPROM
M0 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=885 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=1605 $Y=345 $D=0
M2 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=2535 $Y=345 $D=0
M3 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=885 $Y=2205 $D=16
M4 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1605 $Y=2205 $D=16
M5 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=2535 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKBD1BWP7T I VSS VDD Z
** N=5 EP=4 IP=0 FDC=4
*.SEEDPROM
M0 VSS I 5 VSS N L=1.8e-07 W=4.55e-07 $X=620 $Y=425 $D=0
M1 Z 5 VSS VSS N L=1.8e-07 W=5.2e-07 $X=1440 $Y=360 $D=0
M2 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M3 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1440 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INVD1P5BWP7T I ZN VSS VDD
** N=4 EP=4 IP=0 FDC=4
*.SEEDPROM
M0 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=670 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=5e-07 $X=1440 $Y=345 $D=0
M2 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=670 $Y=2205 $D=16
M3 VDD I ZN VDD P L=1.8e-07 W=6.85e-07 $X=1440 $Y=2890 $D=16
.ENDS
***************************************
.SUBCKT MAOI22D0BWP7T B1 B2 VDD VSS A1 ZN A2
** N=11 EP=7 IP=0 FDC=10
*.SEEDPROM
M0 8 B1 VSS VSS N L=1.8e-07 W=5e-07 $X=460 $Y=845 $D=0
M1 VSS B2 8 VSS N L=1.8e-07 W=5e-07 $X=1180 $Y=845 $D=0
M2 ZN 8 VSS VSS N L=1.8e-07 W=5e-07 $X=1980 $Y=845 $D=0
M3 9 A1 ZN VSS N L=1.8e-07 W=5e-07 $X=2700 $Y=845 $D=0
M4 VSS A2 9 VSS N L=1.8e-07 W=5e-07 $X=3280 $Y=845 $D=0
M5 10 B1 8 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2625 $D=16
M6 VDD B2 10 VDD P L=1.8e-07 W=6.85e-07 $X=1050 $Y=2625 $D=16
M7 11 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1850 $Y=2625 $D=16
M8 ZN A1 11 VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2300 $D=16
M9 11 A2 ZN VDD P L=1.8e-07 W=6.85e-07 $X=3280 $Y=2300 $D=16
.ENDS
***************************************
.SUBCKT OAI31D1BWP7T A1 A2 ZN A3 B VSS VDD
** N=10 EP=7 IP=0 FDC=8
*.SEEDPROM
M0 8 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=680 $Y=345 $D=0
M1 ZN A2 8 VSS N L=1.8e-07 W=1e-06 $X=1400 $Y=345 $D=0
M2 8 A3 ZN VSS N L=1.8e-07 W=1e-06 $X=2160 $Y=345 $D=0
M3 VSS B 8 VSS N L=1.8e-07 W=1e-06 $X=2930 $Y=345 $D=0
M4 9 A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=680 $Y=2205 $D=16
M5 10 A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=1400 $Y=2205 $D=16
M6 ZN A3 10 VDD P L=1.8e-07 W=1.37e-06 $X=2120 $Y=2205 $D=16
M7 VDD B ZN VDD P L=1.8e-07 W=1.37e-06 $X=2930 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OA21D0BWP7T A2 A1 B VDD VSS Z
** N=9 EP=6 IP=0 FDC=8
*.SEEDPROM
M0 7 A2 8 VSS N L=1.8e-07 W=5e-07 $X=460 $Y=750 $D=0
M1 8 A1 7 VSS N L=1.8e-07 W=5e-07 $X=1180 $Y=750 $D=0
M2 VSS B 8 VSS N L=1.8e-07 W=5e-07 $X=1840 $Y=455 $D=0
M3 Z 7 VSS VSS N L=1.8e-07 W=5e-07 $X=2560 $Y=455 $D=0
M4 9 A2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=460 $Y=2350 $D=16
M5 7 A1 9 VDD P L=1.8e-07 W=6.85e-07 $X=1120 $Y=2350 $D=16
M6 VDD B 7 VDD P L=1.8e-07 W=6.85e-07 $X=1840 $Y=2350 $D=16
M7 Z 7 VDD VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2585 $D=16
.ENDS
***************************************
.SUBCKT AOI22D0BWP7T B2 ZN A1 B1 A2 VDD VSS
** N=10 EP=7 IP=0 FDC=8
*.SEEDPROM
M0 8 B2 VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=345 $D=0
M1 ZN B1 8 VSS N L=1.8e-07 W=5e-07 $X=1165 $Y=345 $D=0
M2 9 A1 ZN VSS N L=1.8e-07 W=5e-07 $X=1940 $Y=345 $D=0
M3 VSS A2 9 VSS N L=1.8e-07 W=5e-07 $X=2560 $Y=345 $D=0
M4 10 B2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2755 $D=16
M5 ZN A1 10 VDD P L=1.8e-07 W=6.85e-07 $X=1225 $Y=2555 $D=16
M6 10 A2 ZN VDD P L=1.8e-07 W=6.85e-07 $X=1945 $Y=2555 $D=16
M7 VDD B1 10 VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2890 $D=16
.ENDS
***************************************
.SUBCKT CKND10BWP7T I VDD ZN VSS
** N=4 EP=4 IP=0 FDC=18
*.SEEDPROM
M0 ZN I VSS VSS N L=1.8e-07 W=6.55e-07 $X=1340 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=6.55e-07 $X=2060 $Y=345 $D=0
M2 ZN I VSS VSS N L=1.8e-07 W=6.55e-07 $X=2780 $Y=345 $D=0
M3 VSS I ZN VSS N L=1.8e-07 W=6.55e-07 $X=3500 $Y=345 $D=0
M4 ZN I VSS VSS N L=1.8e-07 W=6.55e-07 $X=4220 $Y=345 $D=0
M5 VSS I ZN VSS N L=1.8e-07 W=6.55e-07 $X=4940 $Y=345 $D=0
M6 ZN I VSS VSS N L=1.8e-07 W=6.55e-07 $X=5660 $Y=345 $D=0
M7 VSS I ZN VSS N L=1.8e-07 W=6.55e-07 $X=6380 $Y=345 $D=0
M8 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M9 VDD I ZN VDD P L=1.8e-07 W=1.565e-06 $X=1340 $Y=2010 $D=16
M10 ZN I VDD VDD P L=1.8e-07 W=1.565e-06 $X=2060 $Y=2010 $D=16
M11 VDD I ZN VDD P L=1.8e-07 W=1.565e-06 $X=2780 $Y=2010 $D=16
M12 ZN I VDD VDD P L=1.8e-07 W=1.565e-06 $X=3500 $Y=2010 $D=16
M13 VDD I ZN VDD P L=1.8e-07 W=1.565e-06 $X=4220 $Y=2010 $D=16
M14 ZN I VDD VDD P L=1.8e-07 W=1.565e-06 $X=4940 $Y=2010 $D=16
M15 VDD I ZN VDD P L=1.8e-07 W=1.565e-06 $X=5660 $Y=2010 $D=16
M16 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=6380 $Y=2205 $D=16
D17 VSS I DN AREA=2.037e-13 PJ=1.81e-06 $X=140 $Y=515 $D=32
.ENDS
***************************************
.SUBCKT ICV_84 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23
+ 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43
+ 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63
+ 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129
** N=425 EP=126 IP=3218 FDC=7873
*.SEEDPROM
M0 422 40 232 4 N L=1.8e-07 W=6.85e-07 $X=227300 $Y=194700 $D=0
M1 4 39 422 4 N L=1.8e-07 W=6.85e-07 $X=227780 $Y=194700 $D=0
M2 237 232 42 4 N L=1.8e-07 W=1e-06 $X=229480 $Y=194545 $D=0
M3 4 31 237 4 N L=1.8e-07 W=1e-06 $X=230200 $Y=194545 $D=0
M4 237 240 4 4 N L=1.8e-07 W=1e-06 $X=230920 $Y=194545 $D=0
M5 44 50 4 4 N L=1.8e-07 W=5e-07 $X=283300 $Y=216875 $D=0
M6 4 50 44 4 N L=1.8e-07 W=5e-07 $X=284020 $Y=216875 $D=0
M7 44 50 4 4 N L=1.8e-07 W=5e-07 $X=284740 $Y=216875 $D=0
M8 4 50 44 4 N L=1.8e-07 W=5e-07 $X=285460 $Y=216875 $D=0
M9 44 54 4 4 N L=1.8e-07 W=5e-07 $X=286180 $Y=216875 $D=0
M10 4 54 44 4 N L=1.8e-07 W=5e-07 $X=286900 $Y=216875 $D=0
M11 44 54 4 4 N L=1.8e-07 W=5e-07 $X=287620 $Y=216875 $D=0
M12 4 54 44 4 N L=1.8e-07 W=5e-07 $X=288340 $Y=216875 $D=0
M13 44 281 4 4 N L=1.8e-07 W=5e-07 $X=289780 $Y=216875 $D=0
M14 4 281 44 4 N L=1.8e-07 W=5e-07 $X=290500 $Y=216875 $D=0
M15 44 281 4 4 N L=1.8e-07 W=5e-07 $X=291220 $Y=216875 $D=0
M16 4 281 44 4 N L=1.8e-07 W=5e-07 $X=291940 $Y=216875 $D=0
M17 4 65 293 4 N L=1.8e-07 W=5.9e-07 $X=296900 $Y=240305 $D=0
M18 293 65 4 4 N L=1.8e-07 W=5.9e-07 $X=297620 $Y=240305 $D=0
M19 4 65 293 4 N L=1.8e-07 W=5.9e-07 $X=298340 $Y=240305 $D=0
M20 293 65 4 4 N L=1.8e-07 W=5.9e-07 $X=299060 $Y=240305 $D=0
M21 4 65 293 4 N L=1.8e-07 W=5.9e-07 $X=299790 $Y=240305 $D=0
M22 68 293 4 4 N L=1.8e-07 W=7.3e-07 $X=300510 $Y=240165 $D=0
M23 4 293 68 4 N L=1.8e-07 W=7.3e-07 $X=301230 $Y=240165 $D=0
M24 68 293 4 4 N L=1.8e-07 W=7.3e-07 $X=301950 $Y=240165 $D=0
M25 4 293 68 4 N L=1.8e-07 W=7.3e-07 $X=302670 $Y=240165 $D=0
M26 68 293 4 4 N L=1.8e-07 W=7.35e-07 $X=304120 $Y=240160 $D=0
M27 4 293 68 4 N L=1.8e-07 W=7.35e-07 $X=304840 $Y=240160 $D=0
M28 68 293 4 4 N L=1.8e-07 W=7.35e-07 $X=305560 $Y=240160 $D=0
M29 4 293 68 4 N L=1.8e-07 W=7.35e-07 $X=306280 $Y=240160 $D=0
M30 68 293 4 4 N L=1.8e-07 W=7.35e-07 $X=307000 $Y=240160 $D=0
M31 423 73 308 4 N L=1.8e-07 W=5e-07 $X=333700 $Y=216540 $D=0
M32 4 74 423 4 N L=1.8e-07 W=5e-07 $X=334200 $Y=216540 $D=0
M33 308 31 4 4 N L=1.8e-07 W=5e-07 $X=334920 $Y=216540 $D=0
M34 4 75 308 4 N L=1.8e-07 W=5e-07 $X=335640 $Y=216540 $D=0
M35 232 40 5 5 P L=1.8e-07 W=6.85e-07 $X=227300 $Y=197020 $D=16
M36 5 39 232 5 P L=1.8e-07 W=6.85e-07 $X=228020 $Y=197020 $D=16
M37 5 232 42 5 P L=1.8e-07 W=1.37e-06 $X=229480 $Y=196405 $D=16
M38 424 31 5 5 P L=1.8e-07 W=1.37e-06 $X=230200 $Y=196405 $D=16
M39 42 240 424 5 P L=1.8e-07 W=1.37e-06 $X=230800 $Y=196405 $D=16
M40 5 50 282 5 P L=1.8e-07 W=1.37e-06 $X=283300 $Y=214145 $D=16
M41 282 50 5 5 P L=1.8e-07 W=1.37e-06 $X=284020 $Y=214145 $D=16
M42 5 50 282 5 P L=1.8e-07 W=1.37e-06 $X=284740 $Y=214145 $D=16
M43 282 50 5 5 P L=1.8e-07 W=1.37e-06 $X=285460 $Y=214145 $D=16
M44 283 54 282 5 P L=1.8e-07 W=1.37e-06 $X=286180 $Y=214145 $D=16
M45 282 54 283 5 P L=1.8e-07 W=1.37e-06 $X=286900 $Y=214145 $D=16
M46 283 54 282 5 P L=1.8e-07 W=1.37e-06 $X=287620 $Y=214145 $D=16
M47 282 54 283 5 P L=1.8e-07 W=1.37e-06 $X=288340 $Y=214145 $D=16
M48 283 281 44 5 P L=1.8e-07 W=1.37e-06 $X=289780 $Y=214145 $D=16
M49 44 281 283 5 P L=1.8e-07 W=1.37e-06 $X=290500 $Y=214145 $D=16
M50 283 281 44 5 P L=1.8e-07 W=1.37e-06 $X=291220 $Y=214145 $D=16
M51 44 281 283 5 P L=1.8e-07 W=1.37e-06 $X=291940 $Y=214145 $D=16
M52 293 65 5 5 P L=1.8e-07 W=1.35e-06 $X=296180 $Y=237665 $D=16
M53 5 65 293 5 P L=1.8e-07 W=1.35e-06 $X=296900 $Y=237665 $D=16
M54 293 65 5 5 P L=1.8e-07 W=1.35e-06 $X=297620 $Y=237665 $D=16
M55 5 65 293 5 P L=1.8e-07 W=1.35e-06 $X=298340 $Y=237665 $D=16
M56 293 65 5 5 P L=1.8e-07 W=1.35e-06 $X=299060 $Y=237665 $D=16
M57 5 65 293 5 P L=1.8e-07 W=1.35e-06 $X=299790 $Y=237665 $D=16
M58 68 293 5 5 P L=1.8e-07 W=1.525e-06 $X=300510 $Y=237665 $D=16
M59 5 293 68 5 P L=1.8e-07 W=1.525e-06 $X=301240 $Y=237665 $D=16
M60 68 293 5 5 P L=1.8e-07 W=1.525e-06 $X=301960 $Y=237665 $D=16
M61 5 293 68 5 P L=1.8e-07 W=1.525e-06 $X=302680 $Y=237665 $D=16
M62 68 293 5 5 P L=1.8e-07 W=1.525e-06 $X=303400 $Y=237665 $D=16
M63 5 293 68 5 P L=1.8e-07 W=1.525e-06 $X=304120 $Y=237665 $D=16
M64 68 293 5 5 P L=1.8e-07 W=1.525e-06 $X=304840 $Y=237665 $D=16
M65 5 293 68 5 P L=1.8e-07 W=1.525e-06 $X=305560 $Y=237665 $D=16
M66 68 293 5 5 P L=1.8e-07 W=1.525e-06 $X=306280 $Y=237665 $D=16
M67 5 293 68 5 P L=1.8e-07 W=1.335e-06 $X=307000 $Y=237665 $D=16
M68 308 73 331 5 P L=1.8e-07 W=1.37e-06 $X=333700 $Y=214145 $D=16
M69 331 74 308 5 P L=1.8e-07 W=1.37e-06 $X=334430 $Y=214145 $D=16
M70 425 31 331 5 P L=1.8e-07 W=1.37e-06 $X=335160 $Y=214145 $D=16
M71 5 75 425 5 P L=1.8e-07 W=1.37e-06 $X=335640 $Y=214145 $D=16
D72 4 65 DN AREA=2.037e-13 PJ=1.81e-06 $X=295700 $Y=240305 $D=32
X255 5 4 DCAPBWP7T $T=156120 155000 0 0 $X=155830 $Y=154765
X256 5 4 DCAPBWP7T $T=156120 233400 1 0 $X=155830 $Y=229190
X257 5 4 DCAPBWP7T $T=163400 225560 0 0 $X=163110 $Y=225325
X258 5 4 DCAPBWP7T $T=184120 241240 1 0 $X=183830 $Y=237030
X259 5 4 DCAPBWP7T $T=185800 186360 0 0 $X=185510 $Y=186125
X260 5 4 DCAPBWP7T $T=186360 202040 1 0 $X=186070 $Y=197830
X261 5 4 DCAPBWP7T $T=195320 162840 1 0 $X=195030 $Y=158630
X262 5 4 DCAPBWP7T $T=195320 194200 1 0 $X=195030 $Y=189990
X263 5 4 DCAPBWP7T $T=195320 202040 1 0 $X=195030 $Y=197830
X264 5 4 DCAPBWP7T $T=195320 209880 1 0 $X=195030 $Y=205670
X265 5 4 DCAPBWP7T $T=195320 241240 1 0 $X=195030 $Y=237030
X266 5 4 DCAPBWP7T $T=198120 186360 0 0 $X=197830 $Y=186125
X267 5 4 DCAPBWP7T $T=209320 194200 1 0 $X=209030 $Y=189990
X268 5 4 DCAPBWP7T $T=209320 209880 1 0 $X=209030 $Y=205670
X269 5 4 DCAPBWP7T $T=222200 162840 1 0 $X=221910 $Y=158630
X270 5 4 DCAPBWP7T $T=222760 209880 0 0 $X=222470 $Y=209645
X271 5 4 DCAPBWP7T $T=240120 194200 0 0 $X=239830 $Y=193965
X272 5 4 DCAPBWP7T $T=240120 225560 1 0 $X=239830 $Y=221350
X273 5 4 DCAPBWP7T $T=258600 170680 0 0 $X=258310 $Y=170445
X274 5 4 DCAPBWP7T $T=260280 209880 0 0 $X=259990 $Y=209645
X275 5 4 DCAPBWP7T $T=279320 162840 1 0 $X=279030 $Y=158630
X276 5 4 DCAPBWP7T $T=321320 186360 1 0 $X=321030 $Y=182150
X277 5 4 DCAPBWP7T $T=321320 202040 1 0 $X=321030 $Y=197830
X278 5 4 DCAPBWP7T $T=321320 217720 1 0 $X=321030 $Y=213510
X279 5 4 DCAPBWP7T $T=333080 225560 0 0 $X=332790 $Y=225325
X280 5 4 DCAPBWP7T $T=335320 186360 1 0 $X=335030 $Y=182150
X281 5 4 DCAPBWP7T $T=339800 233400 0 0 $X=339510 $Y=233165
X282 5 4 DCAPBWP7T $T=363320 162840 0 0 $X=363030 $Y=162605
X283 5 4 DCAPBWP7T $T=363320 202040 1 0 $X=363030 $Y=197830
X284 5 4 DCAPBWP7T $T=363320 209880 1 0 $X=363030 $Y=205670
X285 5 4 DCAPBWP7T $T=363320 209880 0 0 $X=363030 $Y=209645
X286 5 4 DCAPBWP7T $T=372840 202040 1 0 $X=372550 $Y=197830
X287 5 4 DCAPBWP7T $T=372840 209880 0 0 $X=372550 $Y=209645
X288 5 4 DCAPBWP7T $T=375640 202040 0 0 $X=375350 $Y=201805
X289 5 4 DCAPBWP7T $T=377320 241240 1 0 $X=377030 $Y=237030
X290 5 4 DCAPBWP7T $T=386280 178520 0 0 $X=385990 $Y=178285
X291 5 4 DCAPBWP7T $T=386280 186360 0 0 $X=385990 $Y=186125
X292 5 4 DCAPBWP7T $T=405320 155000 0 0 $X=405030 $Y=154765
X293 5 4 DCAPBWP7T $T=405320 170680 1 0 $X=405030 $Y=166470
X294 5 4 DCAPBWP7T $T=405320 186360 0 0 $X=405030 $Y=186125
X295 5 4 DCAPBWP7T $T=405320 209880 1 0 $X=405030 $Y=205670
X296 5 4 DCAPBWP7T $T=405320 225560 0 0 $X=405030 $Y=225325
X297 5 4 DCAPBWP7T $T=405320 241240 1 0 $X=405030 $Y=237030
X298 5 4 DCAPBWP7T $T=414280 170680 0 0 $X=413990 $Y=170445
X299 5 4 DCAPBWP7T $T=414840 202040 1 0 $X=414550 $Y=197830
X300 5 4 DCAPBWP7T $T=415960 186360 1 0 $X=415670 $Y=182150
X301 5 4 DCAPBWP7T $T=421000 170680 0 0 $X=420710 $Y=170445
X302 5 4 DCAPBWP7T $T=427160 202040 1 0 $X=426870 $Y=197830
X303 5 4 DCAPBWP7T $T=432200 225560 0 0 $X=431910 $Y=225325
X304 5 4 DCAPBWP7T $T=439480 202040 1 0 $X=439190 $Y=197830
X305 5 4 DCAPBWP7T $T=440040 217720 0 0 $X=439750 $Y=217485
X306 5 4 DCAPBWP7T $T=447320 209880 0 0 $X=447030 $Y=209645
X307 5 4 DCAPBWP7T $T=447320 225560 1 0 $X=447030 $Y=221350
X308 4 5 DCAP8BWP7T $T=156120 162840 1 0 $X=155830 $Y=158630
X309 4 5 DCAP8BWP7T $T=156120 186360 0 0 $X=155830 $Y=186125
X310 4 5 DCAP8BWP7T $T=156120 241240 1 0 $X=155830 $Y=237030
X311 4 5 DCAP8BWP7T $T=158920 225560 0 0 $X=158630 $Y=225325
X312 4 5 DCAP8BWP7T $T=174040 202040 1 0 $X=173750 $Y=197830
X313 4 5 DCAP8BWP7T $T=177960 155000 0 0 $X=177670 $Y=154765
X314 4 5 DCAP8BWP7T $T=181880 202040 1 0 $X=181590 $Y=197830
X315 4 5 DCAP8BWP7T $T=190840 194200 1 0 $X=190550 $Y=189990
X316 4 5 DCAP8BWP7T $T=190840 202040 1 0 $X=190550 $Y=197830
X317 4 5 DCAP8BWP7T $T=190840 209880 1 0 $X=190550 $Y=205670
X318 4 5 DCAP8BWP7T $T=190840 241240 1 0 $X=190550 $Y=237030
X319 4 5 DCAP8BWP7T $T=191400 225560 0 0 $X=191110 $Y=225325
X320 4 5 DCAP8BWP7T $T=192520 186360 0 0 $X=192230 $Y=186125
X321 4 5 DCAP8BWP7T $T=207080 170680 1 0 $X=206790 $Y=166470
X322 4 5 DCAP8BWP7T $T=207080 225560 0 0 $X=206790 $Y=225325
X323 4 5 DCAP8BWP7T $T=211560 202040 1 0 $X=211270 $Y=197830
X324 4 5 DCAP8BWP7T $T=216040 241240 1 0 $X=215750 $Y=237030
X325 4 5 DCAP8BWP7T $T=218280 186360 0 0 $X=217990 $Y=186125
X326 4 5 DCAP8BWP7T $T=233960 186360 0 0 $X=233670 $Y=186125
X327 4 5 DCAP8BWP7T $T=234520 162840 1 0 $X=234230 $Y=158630
X328 4 5 DCAP8BWP7T $T=234520 209880 0 0 $X=234230 $Y=209645
X329 4 5 DCAP8BWP7T $T=234520 225560 1 0 $X=234230 $Y=221350
X330 4 5 DCAP8BWP7T $T=243480 186360 1 0 $X=243190 $Y=182150
X331 4 5 DCAP8BWP7T $T=249080 186360 0 0 $X=248790 $Y=186125
X332 4 5 DCAP8BWP7T $T=249080 202040 1 0 $X=248790 $Y=197830
X333 4 5 DCAP8BWP7T $T=249080 241240 1 0 $X=248790 $Y=237030
X334 4 5 DCAP8BWP7T $T=267560 170680 0 0 $X=267270 $Y=170445
X335 4 5 DCAP8BWP7T $T=269240 178520 1 0 $X=268950 $Y=174310
X336 4 5 DCAP8BWP7T $T=274280 202040 1 0 $X=273990 $Y=197830
X337 4 5 DCAP8BWP7T $T=274840 162840 1 0 $X=274550 $Y=158630
X338 4 5 DCAP8BWP7T $T=275400 170680 1 0 $X=275110 $Y=166470
X339 4 5 DCAP8BWP7T $T=275400 217720 1 0 $X=275110 $Y=213510
X340 4 5 DCAP8BWP7T $T=275960 170680 0 0 $X=275670 $Y=170445
X341 4 5 DCAP8BWP7T $T=275960 194200 1 0 $X=275670 $Y=189990
X342 4 5 DCAP8BWP7T $T=275960 202040 0 0 $X=275670 $Y=201805
X343 4 5 DCAP8BWP7T $T=275960 217720 0 0 $X=275670 $Y=217485
X344 4 5 DCAP8BWP7T $T=275960 241240 1 0 $X=275670 $Y=237030
X345 4 5 DCAP8BWP7T $T=276520 178520 1 0 $X=276230 $Y=174310
X346 4 5 DCAP8BWP7T $T=276520 225560 0 0 $X=276230 $Y=225325
X347 4 5 DCAP8BWP7T $T=285480 209880 0 0 $X=285190 $Y=209645
X348 4 5 DCAP8BWP7T $T=291080 178520 1 0 $X=290790 $Y=174310
X349 4 5 DCAP8BWP7T $T=291080 241240 1 0 $X=290790 $Y=237030
X350 4 5 DCAP8BWP7T $T=293320 233400 0 0 $X=293030 $Y=233165
X351 4 5 DCAP8BWP7T $T=316840 202040 1 0 $X=316550 $Y=197830
X352 4 5 DCAP8BWP7T $T=316840 217720 1 0 $X=316550 $Y=213510
X353 4 5 DCAP8BWP7T $T=317960 178520 1 0 $X=317670 $Y=174310
X354 4 5 DCAP8BWP7T $T=317960 217720 0 0 $X=317670 $Y=217485
X355 4 5 DCAP8BWP7T $T=317960 241240 1 0 $X=317670 $Y=237030
X356 4 5 DCAP8BWP7T $T=318520 170680 0 0 $X=318230 $Y=170445
X357 4 5 DCAP8BWP7T $T=318520 233400 0 0 $X=318230 $Y=233165
X358 4 5 DCAP8BWP7T $T=326920 202040 1 0 $X=326630 $Y=197830
X359 4 5 DCAP8BWP7T $T=333080 209880 1 0 $X=332790 $Y=205670
X360 4 5 DCAP8BWP7T $T=340360 186360 0 0 $X=340070 $Y=186125
X361 4 5 DCAP8BWP7T $T=351000 155000 0 0 $X=350710 $Y=154765
X362 4 5 DCAP8BWP7T $T=351000 170680 1 0 $X=350710 $Y=166470
X363 4 5 DCAP8BWP7T $T=353240 170680 0 0 $X=352950 $Y=170445
X364 4 5 DCAP8BWP7T $T=358840 202040 1 0 $X=358550 $Y=197830
X365 4 5 DCAP8BWP7T $T=358840 209880 1 0 $X=358550 $Y=205670
X366 4 5 DCAP8BWP7T $T=359960 202040 0 0 $X=359670 $Y=201805
X367 4 5 DCAP8BWP7T $T=360520 155000 0 0 $X=360230 $Y=154765
X368 4 5 DCAP8BWP7T $T=360520 170680 0 0 $X=360230 $Y=170445
X369 4 5 DCAP8BWP7T $T=360520 186360 1 0 $X=360230 $Y=182150
X370 4 5 DCAP8BWP7T $T=360520 225560 0 0 $X=360230 $Y=225325
X371 4 5 DCAP8BWP7T $T=366120 178520 1 0 $X=365830 $Y=174310
X372 4 5 DCAP8BWP7T $T=368360 202040 1 0 $X=368070 $Y=197830
X373 4 5 DCAP8BWP7T $T=368360 209880 0 0 $X=368070 $Y=209645
X374 4 5 DCAP8BWP7T $T=375080 162840 1 0 $X=374790 $Y=158630
X375 4 5 DCAP8BWP7T $T=377320 209880 0 0 $X=377030 $Y=209645
X376 4 5 DCAP8BWP7T $T=381800 186360 0 0 $X=381510 $Y=186125
X377 4 5 DCAP8BWP7T $T=401400 225560 1 0 $X=401110 $Y=221350
X378 4 5 DCAP8BWP7T $T=401960 233400 0 0 $X=401670 $Y=233165
X379 4 5 DCAP8BWP7T $T=402520 162840 1 0 $X=402230 $Y=158630
X380 4 5 DCAP8BWP7T $T=402520 178520 1 0 $X=402230 $Y=174310
X381 4 5 DCAP8BWP7T $T=402520 217720 0 0 $X=402230 $Y=217485
X382 4 5 DCAP8BWP7T $T=408120 178520 0 0 $X=407830 $Y=178285
X383 4 5 DCAP8BWP7T $T=408120 217720 1 0 $X=407830 $Y=213510
X384 4 5 DCAP8BWP7T $T=408120 217720 0 0 $X=407830 $Y=217485
X385 4 5 DCAP8BWP7T $T=412040 209880 0 0 $X=411750 $Y=209645
X386 4 5 DCAP8BWP7T $T=414280 186360 0 0 $X=413990 $Y=186125
X387 4 5 DCAP8BWP7T $T=429400 186360 1 0 $X=429110 $Y=182150
X388 4 5 DCAP8BWP7T $T=435560 178520 1 0 $X=435270 $Y=174310
X389 4 5 DCAP8BWP7T $T=443960 178520 0 0 $X=443670 $Y=178285
X390 4 5 DCAP8BWP7T $T=443960 209880 1 0 $X=443670 $Y=205670
X391 4 5 DCAP8BWP7T $T=444520 155000 0 0 $X=444230 $Y=154765
X392 4 5 DCAP8BWP7T $T=444520 178520 1 0 $X=444230 $Y=174310
X393 4 5 DCAP8BWP7T $T=444520 202040 1 0 $X=444230 $Y=197830
X394 4 5 DCAP8BWP7T $T=444520 217720 0 0 $X=444230 $Y=217485
X395 4 5 DCAP8BWP7T $T=444520 225560 0 0 $X=444230 $Y=225325
X396 4 5 DCAP8BWP7T $T=444520 241240 1 0 $X=444230 $Y=237030
X397 4 5 DCAP4BWP7T $T=156120 162840 0 0 $X=155830 $Y=162605
X398 4 5 DCAP4BWP7T $T=166200 162840 1 0 $X=165910 $Y=158630
X399 4 5 DCAP4BWP7T $T=175160 202040 0 0 $X=174870 $Y=201805
X400 4 5 DCAP4BWP7T $T=176280 194200 1 0 $X=175990 $Y=189990
X401 4 5 DCAP4BWP7T $T=193640 170680 0 0 $X=193350 $Y=170445
X402 4 5 DCAP4BWP7T $T=194200 170680 1 0 $X=193910 $Y=166470
X403 4 5 DCAP4BWP7T $T=194200 178520 0 0 $X=193910 $Y=178285
X404 4 5 DCAP4BWP7T $T=194200 194200 0 0 $X=193910 $Y=193965
X405 4 5 DCAP4BWP7T $T=222200 178520 1 0 $X=221910 $Y=174310
X406 4 5 DCAP4BWP7T $T=235640 155000 0 0 $X=235350 $Y=154765
X407 4 5 DCAP4BWP7T $T=236200 202040 1 0 $X=235910 $Y=197830
X408 4 5 DCAP4BWP7T $T=240120 194200 1 0 $X=239830 $Y=189990
X409 4 5 DCAP4BWP7T $T=240120 202040 0 0 $X=239830 $Y=201805
X410 4 5 DCAP4BWP7T $T=251320 194200 1 0 $X=251030 $Y=189990
X411 4 5 DCAP4BWP7T $T=256920 186360 1 0 $X=256630 $Y=182150
X412 4 5 DCAP4BWP7T $T=278200 155000 0 0 $X=277910 $Y=154765
X413 4 5 DCAP4BWP7T $T=278760 209880 0 0 $X=278470 $Y=209645
X414 4 5 DCAP4BWP7T $T=282120 225560 1 0 $X=281830 $Y=221350
X415 4 5 DCAP4BWP7T $T=284920 202040 1 0 $X=284630 $Y=197830
X416 4 5 DCAP4BWP7T $T=301720 217720 1 0 $X=301430 $Y=213510
X417 4 5 DCAP4BWP7T $T=310120 241240 1 0 $X=309830 $Y=237030
X418 4 5 DCAP4BWP7T $T=320200 225560 1 0 $X=319910 $Y=221350
X419 4 5 DCAP4BWP7T $T=320760 194200 1 0 $X=320470 $Y=189990
X420 4 5 DCAP4BWP7T $T=320760 194200 0 0 $X=320470 $Y=193965
X421 4 5 DCAP4BWP7T $T=320760 202040 0 0 $X=320470 $Y=201805
X422 4 5 DCAP4BWP7T $T=320760 209880 0 0 $X=320470 $Y=209645
X423 4 5 DCAP4BWP7T $T=324120 178520 1 0 $X=323830 $Y=174310
X424 4 5 DCAP4BWP7T $T=361080 209880 0 0 $X=360790 $Y=209645
X425 4 5 DCAP4BWP7T $T=362760 217720 0 0 $X=362470 $Y=217485
X426 4 5 DCAP4BWP7T $T=366120 225560 0 0 $X=365830 $Y=225325
X427 4 5 DCAP4BWP7T $T=366120 233400 1 0 $X=365830 $Y=229190
X428 4 5 DCAP4BWP7T $T=368920 186360 0 0 $X=368630 $Y=186125
X429 4 5 DCAP4BWP7T $T=377880 202040 1 0 $X=377590 $Y=197830
X430 4 5 DCAP4BWP7T $T=384040 178520 0 0 $X=383750 $Y=178285
X431 4 5 DCAP4BWP7T $T=397480 217720 0 0 $X=397190 $Y=217485
X432 4 5 DCAP4BWP7T $T=403080 186360 0 0 $X=402790 $Y=186125
X433 4 5 DCAP4BWP7T $T=404200 209880 0 0 $X=403910 $Y=209645
X434 4 5 DCAP4BWP7T $T=408120 186360 0 0 $X=407830 $Y=186125
X435 4 5 DCAP4BWP7T $T=408120 194200 0 0 $X=407830 $Y=193965
X436 4 5 DCAP4BWP7T $T=408120 225560 0 0 $X=407830 $Y=225325
X437 4 5 DCAP4BWP7T $T=412040 170680 0 0 $X=411750 $Y=170445
X438 4 5 DCAP4BWP7T $T=412600 202040 1 0 $X=412310 $Y=197830
X439 4 5 DCAP4BWP7T $T=429960 225560 0 0 $X=429670 $Y=225325
X440 4 5 DCAP4BWP7T $T=438920 209880 1 0 $X=438630 $Y=205670
X441 4 5 DCAP4BWP7T $T=445640 170680 0 0 $X=445350 $Y=170445
X442 4 5 DCAP4BWP7T $T=445640 186360 0 0 $X=445350 $Y=186125
X443 4 5 DCAP4BWP7T $T=446200 194200 1 0 $X=445910 $Y=189990
X444 4 5 ICV_40 $T=156120 170680 0 0 $X=155830 $Y=170445
X445 4 5 ICV_40 $T=189160 233400 1 0 $X=188870 $Y=229190
X446 4 5 ICV_40 $T=189720 178520 1 0 $X=189430 $Y=174310
X447 4 5 ICV_40 $T=189720 202040 0 0 $X=189430 $Y=201805
X448 4 5 ICV_40 $T=189720 209880 0 0 $X=189430 $Y=209645
X449 4 5 ICV_40 $T=215480 162840 1 0 $X=215190 $Y=158630
X450 4 5 ICV_40 $T=216040 202040 0 0 $X=215750 $Y=201805
X451 4 5 ICV_40 $T=216040 209880 0 0 $X=215750 $Y=209645
X452 4 5 ICV_40 $T=231720 170680 1 0 $X=231430 $Y=166470
X453 4 5 ICV_40 $T=231720 178520 1 0 $X=231430 $Y=174310
X454 4 5 ICV_40 $T=231720 194200 0 0 $X=231430 $Y=193965
X455 4 5 ICV_40 $T=231720 217720 0 0 $X=231430 $Y=217485
X456 4 5 ICV_40 $T=232280 178520 0 0 $X=231990 $Y=178285
X457 4 5 ICV_40 $T=232280 233400 0 0 $X=231990 $Y=233165
X458 4 5 ICV_40 $T=245720 194200 0 0 $X=245430 $Y=193965
X459 4 5 ICV_40 $T=251880 170680 0 0 $X=251590 $Y=170445
X460 4 5 ICV_40 $T=255240 155000 0 0 $X=254950 $Y=154765
X461 4 5 ICV_40 $T=263640 225560 1 0 $X=263350 $Y=221350
X462 4 5 ICV_40 $T=264760 209880 0 0 $X=264470 $Y=209645
X463 4 5 ICV_40 $T=273160 186360 1 0 $X=272870 $Y=182150
X464 4 5 ICV_40 $T=273160 225560 1 0 $X=272870 $Y=221350
X465 4 5 ICV_40 $T=273720 186360 0 0 $X=273430 $Y=186125
X466 4 5 ICV_40 $T=274280 194200 0 0 $X=273990 $Y=193965
X467 4 5 ICV_40 $T=316280 162840 1 0 $X=315990 $Y=158630
X468 4 5 ICV_40 $T=316280 186360 0 0 $X=315990 $Y=186125
X469 4 5 ICV_40 $T=333080 170680 0 0 $X=332790 $Y=170445
X470 4 5 ICV_40 $T=333080 233400 0 0 $X=332790 $Y=233165
X471 4 5 ICV_40 $T=333080 241240 1 0 $X=332790 $Y=237030
X472 4 5 ICV_40 $T=357720 186360 0 0 $X=357430 $Y=186125
X473 4 5 ICV_40 $T=358280 217720 1 0 $X=357990 $Y=213510
X474 4 5 ICV_40 $T=368920 202040 0 0 $X=368630 $Y=201805
X475 4 5 ICV_40 $T=368920 217720 1 0 $X=368630 $Y=213510
X476 4 5 ICV_40 $T=371720 225560 0 0 $X=371430 $Y=225325
X477 4 5 ICV_40 $T=375080 225560 1 0 $X=374790 $Y=221350
X478 4 5 ICV_40 $T=398600 225560 0 0 $X=398310 $Y=225325
X479 4 5 ICV_40 $T=398600 241240 1 0 $X=398310 $Y=237030
X480 4 5 ICV_40 $T=399720 178520 0 0 $X=399430 $Y=178285
X481 4 5 ICV_40 $T=399720 202040 1 0 $X=399430 $Y=197830
X482 4 5 ICV_40 $T=400280 194200 0 0 $X=399990 $Y=193965
X483 4 5 ICV_40 $T=400280 233400 1 0 $X=399990 $Y=229190
X484 4 5 ICV_40 $T=415960 178520 0 0 $X=415670 $Y=178285
X485 4 5 ICV_40 $T=424920 217720 1 0 $X=424630 $Y=213510
X486 4 5 ICV_40 $T=426040 155000 0 0 $X=425750 $Y=154765
X487 4 5 ICV_40 $T=441160 194200 0 0 $X=440870 $Y=193965
X488 4 5 ICV_40 $T=442280 217720 1 0 $X=441990 $Y=213510
X489 7 5 139 6 4 NR2D1BWP7T $T=156120 178520 1 0 $X=155830 $Y=174310
X490 7 5 135 133 4 NR2D1BWP7T $T=158360 178520 1 180 $X=155830 $Y=178285
X491 8 5 136 6 4 NR2D1BWP7T $T=158360 194200 0 180 $X=155830 $Y=189990
X492 133 5 142 14 4 NR2D1BWP7T $T=156120 194200 0 0 $X=155830 $Y=193965
X493 8 5 137 133 4 NR2D1BWP7T $T=158360 202040 1 180 $X=155830 $Y=201805
X494 134 5 11 9 4 NR2D1BWP7T $T=160040 155000 1 180 $X=157510 $Y=154765
X495 15 5 13 9 4 NR2D1BWP7T $T=160040 233400 0 180 $X=157510 $Y=229190
X496 134 5 146 133 4 NR2D1BWP7T $T=159480 162840 0 0 $X=159190 $Y=162605
X497 16 5 145 14 4 NR2D1BWP7T $T=162280 233400 0 180 $X=159750 $Y=229190
X498 133 5 151 15 4 NR2D1BWP7T $T=161720 241240 1 0 $X=161430 $Y=237030
X499 134 5 155 21 4 NR2D1BWP7T $T=175160 162840 1 0 $X=174870 $Y=158630
X500 16 5 164 15 4 NR2D1BWP7T $T=177400 241240 0 180 $X=174870 $Y=237030
X501 134 5 143 6 4 NR2D1BWP7T $T=177400 186360 0 0 $X=177110 $Y=186125
X502 14 5 167 6 4 NR2D1BWP7T $T=177400 241240 1 0 $X=177110 $Y=237030
X503 7 5 182 22 4 NR2D1BWP7T $T=189720 202040 1 180 $X=187190 $Y=201805
X504 16 5 171 7 4 NR2D1BWP7T $T=189720 209880 1 180 $X=187190 $Y=209645
X505 8 5 187 21 4 NR2D1BWP7T $T=188600 241240 1 0 $X=188310 $Y=237030
X506 203 5 201 9 4 NR2D1BWP7T $T=208760 217720 0 180 $X=206230 $Y=213510
X507 134 5 220 16 4 NR2D1BWP7T $T=224440 209880 0 0 $X=224150 $Y=209645
X508 31 5 244 242 4 NR2D1BWP7T $T=240680 170680 0 0 $X=240390 $Y=170445
X509 251 5 253 257 4 NR2D1BWP7T $T=253560 202040 1 0 $X=253270 $Y=197830
X510 16 5 205 8 4 NR2D1BWP7T $T=261400 225560 1 180 $X=258870 $Y=225325
X511 203 5 270 257 4 NR2D1BWP7T $T=272040 209880 0 0 $X=271750 $Y=209645
X512 54 5 272 277 4 NR2D1BWP7T $T=282680 194200 1 0 $X=282390 $Y=189990
X513 203 5 284 277 4 NR2D1BWP7T $T=282680 194200 0 0 $X=282390 $Y=193965
X514 281 5 239 203 4 NR2D1BWP7T $T=285480 209880 1 180 $X=282950 $Y=209645
X515 203 5 265 255 4 NR2D1BWP7T $T=287720 225560 0 180 $X=285190 $Y=221350
X516 281 5 287 62 4 NR2D1BWP7T $T=293880 202040 0 180 $X=291350 $Y=197830
X517 281 5 289 290 4 NR2D1BWP7T $T=293880 202040 1 0 $X=293590 $Y=197830
X518 281 5 298 67 4 NR2D1BWP7T $T=300040 225560 1 0 $X=299750 $Y=221350
X519 251 5 302 277 4 NR2D1BWP7T $T=300600 202040 1 0 $X=300310 $Y=197830
X520 281 5 312 70 4 NR2D1BWP7T $T=312920 241240 1 0 $X=312630 $Y=237030
X521 62 5 321 257 4 NR2D1BWP7T $T=315720 225560 0 0 $X=315430 $Y=225325
X522 290 5 71 9 4 NR2D1BWP7T $T=317960 241240 0 180 $X=315430 $Y=237030
X523 281 5 267 251 4 NR2D1BWP7T $T=326920 202040 0 180 $X=324390 $Y=197830
X524 277 5 292 62 4 NR2D1BWP7T $T=326920 217720 0 180 $X=324390 $Y=213510
X525 277 5 322 290 4 NR2D1BWP7T $T=324680 217720 0 0 $X=324390 $Y=217485
X526 251 5 323 324 4 NR2D1BWP7T $T=326920 202040 0 0 $X=326630 $Y=201805
X527 54 5 294 257 4 NR2D1BWP7T $T=337000 186360 1 0 $X=336710 $Y=182150
X528 203 5 306 324 4 NR2D1BWP7T $T=340360 186360 1 180 $X=337830 $Y=186125
X529 54 5 311 324 4 NR2D1BWP7T $T=338680 209880 1 0 $X=338390 $Y=205670
X530 67 5 343 255 4 NR2D1BWP7T $T=368920 194200 1 180 $X=366390 $Y=193965
X531 91 5 88 9 4 NR2D1BWP7T $T=370040 233400 1 180 $X=367510 $Y=233165
X532 5 4 DCAP64BWP7T $T=158360 178520 0 0 $X=158070 $Y=178285
X533 5 4 DCAP64BWP7T $T=284920 194200 1 0 $X=284630 $Y=189990
X534 5 4 DCAP64BWP7T $T=284920 202040 0 0 $X=284630 $Y=201805
X535 5 4 DCAP64BWP7T $T=285480 186360 1 0 $X=285190 $Y=182150
X536 5 4 DCAP64BWP7T $T=327480 162840 0 0 $X=327190 $Y=162605
X537 5 4 DCAP64BWP7T $T=411480 225560 1 0 $X=411190 $Y=221350
X538 4 5 ICV_46 $T=408120 162840 0 0 $X=407830 $Y=162605
X539 4 5 ICV_46 $T=408120 170680 1 0 $X=407830 $Y=166470
X540 4 5 ICV_46 $T=408120 233400 0 0 $X=407830 $Y=233165
X587 4 5 ICV_47 $T=156120 186360 1 0 $X=155830 $Y=182150
X588 4 5 ICV_47 $T=156120 217720 0 0 $X=155830 $Y=217485
X589 4 5 ICV_47 $T=156120 225560 1 0 $X=155830 $Y=221350
X590 4 5 ICV_47 $T=156120 233400 0 0 $X=155830 $Y=233165
X591 4 5 ICV_47 $T=198120 186360 1 0 $X=197830 $Y=182150
X592 4 5 ICV_47 $T=240120 162840 0 0 $X=239830 $Y=162605
X593 4 5 ICV_47 $T=240120 178520 0 0 $X=239830 $Y=178285
X594 4 5 ICV_47 $T=240120 233400 1 0 $X=239830 $Y=229190
X595 4 5 ICV_47 $T=282120 155000 0 0 $X=281830 $Y=154765
X596 4 5 ICV_47 $T=282120 170680 1 0 $X=281830 $Y=166470
X597 4 5 ICV_47 $T=282120 178520 0 0 $X=281830 $Y=178285
X598 4 5 ICV_47 $T=282120 209880 1 0 $X=281830 $Y=205670
X599 4 5 ICV_47 $T=324120 178520 0 0 $X=323830 $Y=178285
X600 4 5 ICV_47 $T=324120 194200 1 0 $X=323830 $Y=189990
X601 4 5 ICV_47 $T=324120 194200 0 0 $X=323830 $Y=193965
X602 4 5 ICV_47 $T=324120 225560 1 0 $X=323830 $Y=221350
X603 4 5 ICV_47 $T=366120 194200 1 0 $X=365830 $Y=189990
X604 5 4 DCAP32BWP7T $T=156120 202040 1 0 $X=155830 $Y=197830
X605 5 4 DCAP32BWP7T $T=156120 209880 1 0 $X=155830 $Y=205670
X606 5 4 DCAP32BWP7T $T=156120 209880 0 0 $X=155830 $Y=209645
X607 5 4 DCAP32BWP7T $T=158360 194200 1 0 $X=158070 $Y=189990
X608 5 4 DCAP32BWP7T $T=161720 162840 0 0 $X=161430 $Y=162605
X609 5 4 DCAP32BWP7T $T=198120 202040 0 0 $X=197830 $Y=201805
X610 5 4 DCAP32BWP7T $T=198120 209880 0 0 $X=197830 $Y=209645
X611 5 4 DCAP32BWP7T $T=198120 241240 1 0 $X=197830 $Y=237030
X612 5 4 DCAP32BWP7T $T=208760 217720 1 0 $X=208470 $Y=213510
X613 5 4 DCAP32BWP7T $T=211560 233400 1 0 $X=211270 $Y=229190
X614 5 4 DCAP32BWP7T $T=217720 155000 0 0 $X=217430 $Y=154765
X615 5 4 DCAP32BWP7T $T=218280 202040 1 0 $X=217990 $Y=197830
X616 5 4 DCAP32BWP7T $T=220520 194200 1 0 $X=220230 $Y=189990
X617 5 4 DCAP32BWP7T $T=240120 217720 1 0 $X=239830 $Y=213510
X618 5 4 DCAP32BWP7T $T=253560 233400 0 0 $X=253270 $Y=233165
X619 5 4 DCAP32BWP7T $T=255800 186360 0 0 $X=255510 $Y=186125
X620 5 4 DCAP32BWP7T $T=263080 209880 1 0 $X=262790 $Y=205670
X621 5 4 DCAP32BWP7T $T=282120 225560 0 0 $X=281830 $Y=225325
X622 5 4 DCAP32BWP7T $T=300600 233400 0 0 $X=300310 $Y=233165
X623 5 4 DCAP32BWP7T $T=302280 225560 1 0 $X=301990 $Y=221350
X624 5 4 DCAP32BWP7T $T=302840 209880 0 0 $X=302550 $Y=209645
X625 5 4 DCAP32BWP7T $T=324120 155000 0 0 $X=323830 $Y=154765
X626 5 4 DCAP32BWP7T $T=324120 170680 1 0 $X=323830 $Y=166470
X627 5 4 DCAP32BWP7T $T=337560 233400 1 0 $X=337270 $Y=229190
X628 5 4 DCAP32BWP7T $T=340920 209880 1 0 $X=340630 $Y=205670
X629 5 4 DCAP32BWP7T $T=342600 186360 1 0 $X=342310 $Y=182150
X630 5 4 DCAP32BWP7T $T=343160 209880 0 0 $X=342870 $Y=209645
X631 5 4 DCAP32BWP7T $T=366120 178520 0 0 $X=365830 $Y=178285
X632 5 4 DCAP32BWP7T $T=373400 233400 1 0 $X=373110 $Y=229190
X633 5 4 DCAP32BWP7T $T=377880 162840 0 0 $X=377590 $Y=162605
X634 5 4 DCAP32BWP7T $T=381800 186360 1 0 $X=381510 $Y=182150
X635 5 4 DCAP32BWP7T $T=408120 155000 0 0 $X=407830 $Y=154765
X636 5 4 DCAP32BWP7T $T=408120 194200 1 0 $X=407830 $Y=189990
X637 5 4 DCAP32BWP7T $T=408120 202040 0 0 $X=407830 $Y=201805
X638 5 4 DCAP32BWP7T $T=408120 233400 1 0 $X=407830 $Y=229190
X639 5 4 DCAP32BWP7T $T=426040 178520 0 0 $X=425750 $Y=178285
X640 5 4 DCAP32BWP7T $T=429400 209880 0 0 $X=429110 $Y=209645
X641 5 4 DCAP32BWP7T $T=429960 233400 1 0 $X=429670 $Y=229190
X642 135 145 143 140 5 4 132 FA1D0BWP7T $T=169000 217720 0 180 $X=155830 $Y=213510
X643 147 140 158 161 5 4 152 FA1D0BWP7T $T=161720 186360 0 0 $X=161430 $Y=186125
X644 150 132 159 160 5 4 163 FA1D0BWP7T $T=162280 202040 0 0 $X=161990 $Y=201805
X645 152 154 160 162 5 4 165 FA1D0BWP7T $T=162840 170680 0 0 $X=162550 $Y=170445
X646 164 137 155 150 5 4 18 FA1D0BWP7T $T=177960 225560 1 180 $X=164790 $Y=225325
X647 175 166 139 159 5 4 156 FA1D0BWP7T $T=183000 217720 0 180 $X=169830 $Y=213510
X648 153 173 179 181 5 4 184 FA1D0BWP7T $T=176840 178520 1 0 $X=176550 $Y=174310
X649 138 136 142 186 5 4 191 FA1D0BWP7T $T=178520 225560 0 0 $X=178230 $Y=225325
X650 168 182 205 207 5 4 183 FA1D0BWP7T $T=198680 202040 1 0 $X=198390 $Y=197830
X651 29 186 156 198 5 4 211 FA1D0BWP7T $T=198680 233400 1 0 $X=198390 $Y=229190
X652 210 191 223 224 5 4 225 FA1D0BWP7T $T=209880 217720 0 0 $X=209590 $Y=217485
X653 167 151 187 210 5 4 37 FA1D0BWP7T $T=210440 233400 0 0 $X=210150 $Y=233165
X654 216 228 211 231 5 4 241 FA1D0BWP7T $T=221640 225560 1 0 $X=221350 $Y=221350
X655 193 38 43 223 5 4 45 FA1D0BWP7T $T=221640 241240 1 0 $X=221350 $Y=237030
X656 51 224 49 228 5 4 46 FA1D0BWP7T $T=253560 233400 1 180 $X=240390 $Y=233165
X657 274 233 261 242 5 4 217 FA1D0BWP7T $T=273160 186360 0 180 $X=259990 $Y=182150
X658 180 265 267 269 5 4 273 FA1D0BWP7T $T=261400 202040 1 0 $X=261110 $Y=197830
X659 285 286 275 264 5 4 279 FA1D0BWP7T $T=296120 170680 1 180 $X=282950 $Y=170445
X660 284 287 294 286 5 4 300 FA1D0BWP7T $T=289400 186360 0 0 $X=289110 $Y=186125
X661 250 253 292 297 5 4 301 FA1D0BWP7T $T=289960 209880 0 0 $X=289670 $Y=209645
X662 279 266 304 291 5 4 314 FA1D0BWP7T $T=296120 178520 1 0 $X=295830 $Y=174310
X663 271 254 270 305 5 4 318 FA1D0BWP7T $T=303400 186360 0 0 $X=303110 $Y=186125
X664 289 302 311 316 5 4 319 FA1D0BWP7T $T=303960 202040 1 0 $X=303670 $Y=197830
X665 298 306 313 317 5 4 320 FA1D0BWP7T $T=303960 217720 1 0 $X=303670 $Y=213510
X666 316 300 305 304 5 4 303 FA1D0BWP7T $T=318520 170680 1 180 $X=305350 $Y=170445
X667 317 326 319 329 5 4 336 FA1D0BWP7T $T=324680 186360 0 0 $X=324390 $Y=186125
X668 321 322 323 335 5 4 337 FA1D0BWP7T $T=324680 233400 1 0 $X=324390 $Y=229190
X669 297 329 318 310 5 4 338 FA1D0BWP7T $T=326360 178520 1 0 $X=326070 $Y=174310
X670 330 333 338 346 5 4 347 FA1D0BWP7T $T=331400 162840 1 0 $X=331110 $Y=158630
X671 295 320 339 348 5 4 77 FA1D0BWP7T $T=332520 202040 1 0 $X=332230 $Y=197830
X672 334 301 335 350 5 4 78 FA1D0BWP7T $T=334760 225560 0 0 $X=334470 $Y=225325
X673 350 348 336 333 5 4 341 FA1D0BWP7T $T=353240 170680 1 180 $X=340070 $Y=170445
X674 362 312 353 334 5 4 79 FA1D0BWP7T $T=360520 225560 1 180 $X=347350 $Y=225325
X675 10 4 5 134 INVD1BWP7T $T=158360 170680 0 180 $X=156390 $Y=166470
X676 20 4 5 133 INVD1BWP7T $T=165640 241240 0 180 $X=163670 $Y=237030
X677 157 4 5 19 INVD1BWP7T $T=171240 162840 0 180 $X=169270 $Y=158630
X678 189 4 5 7 INVD1BWP7T $T=200360 217720 0 180 $X=198390 $Y=213510
X679 195 4 5 190 INVD1BWP7T $T=201480 162840 1 0 $X=201190 $Y=158630
X680 197 4 5 27 INVD1BWP7T $T=203160 162840 1 0 $X=202870 $Y=158630
X681 200 4 5 30 INVD1BWP7T $T=204840 162840 1 0 $X=204550 $Y=158630
X682 212 4 5 208 INVD1BWP7T $T=212120 155000 1 180 $X=210150 $Y=154765
X683 61 4 5 277 INVD1BWP7T $T=274840 225560 0 0 $X=274550 $Y=225325
X684 280 4 5 62 INVD1BWP7T $T=300040 225560 0 180 $X=298070 $Y=221350
X685 72 4 5 257 INVD1BWP7T $T=329160 217720 1 0 $X=328870 $Y=213510
X686 307 4 5 209 INVD1BWP7T $T=349320 162840 1 0 $X=349030 $Y=158630
X687 356 4 5 67 INVD1BWP7T $T=355480 162840 0 180 $X=353510 $Y=158630
X688 364 4 5 290 INVD1BWP7T $T=368360 202040 0 180 $X=366390 $Y=197830
X689 141 4 5 138 CKBD0BWP7T $T=158920 225560 1 180 $X=156390 $Y=225325
X788 148 4 144 12 5 ND2D1BWP7T $T=160600 202040 1 180 $X=158070 $Y=201805
X789 238 4 235 41 5 ND2D1BWP7T $T=231720 178520 0 180 $X=229190 $Y=174310
X790 52 4 194 41 5 ND2D1BWP7T $T=253560 186360 0 0 $X=253270 $Y=186125
X791 189 4 59 60 5 ND2D1BWP7T $T=271480 241240 1 0 $X=271190 $Y=237030
X792 280 4 252 41 5 ND2D1BWP7T $T=284920 186360 1 180 $X=282390 $Y=186125
X793 10 4 170 55 5 ND2D1BWP7T $T=284920 202040 1 180 $X=282390 $Y=201805
X794 148 4 196 55 5 ND2D1BWP7T $T=329160 217720 0 180 $X=326630 $Y=213510
X795 280 4 328 76 5 ND2D1BWP7T $T=339240 209880 1 180 $X=336710 $Y=209645
X796 364 4 360 41 5 ND2D1BWP7T $T=368920 186360 1 180 $X=366390 $Y=186125
X797 92 4 357 238 5 ND2D1BWP7T $T=368920 202040 1 180 $X=366390 $Y=201805
X798 41 4 351 89 5 ND2D1BWP7T $T=368920 217720 0 180 $X=366390 $Y=213510
X799 93 4 358 52 5 ND2D1BWP7T $T=370600 233400 0 180 $X=368070 $Y=229190
X800 349 4 340 94 5 ND2D1BWP7T $T=369480 225560 0 0 $X=369190 $Y=225325
X817 149 4 5 147 INVD0BWP7T $T=163400 162840 0 180 $X=161430 $Y=158630
X818 176 4 5 154 INVD0BWP7T $T=181320 186360 1 180 $X=179350 $Y=186125
X819 184 4 5 188 INVD0BWP7T $T=201480 162840 0 180 $X=199510 $Y=158630
X820 214 4 5 174 INVD0BWP7T $T=212680 178520 1 180 $X=210710 $Y=178285
X821 207 4 5 179 INVD0BWP7T $T=218280 202040 0 180 $X=216310 $Y=197830
X822 264 4 5 259 INVD0BWP7T $T=264760 155000 1 180 $X=262790 $Y=154765
X823 249 4 5 256 INVD0BWP7T $T=267560 155000 0 0 $X=267270 $Y=154765
X824 273 4 5 260 INVD0BWP7T $T=275400 170680 0 180 $X=273430 $Y=166470
X825 269 4 5 261 INVD0BWP7T $T=282680 162840 1 0 $X=282390 $Y=158630
X826 276 4 5 285 INVD0BWP7T $T=289400 162840 1 0 $X=289110 $Y=158630
X827 325 4 5 330 INVD0BWP7T $T=347640 162840 1 0 $X=347350 $Y=158630
X828 76 4 5 324 INVD0BWP7T $T=368360 209880 1 180 $X=366390 $Y=209645
X829 146 153 17 149 4 5 OAI21D0BWP7T $T=163400 162840 1 0 $X=163110 $Y=158630
X830 163 199 198 165 4 5 OAI21D0BWP7T $T=206520 217720 0 180 $X=203430 $Y=213510
X831 219 218 217 34 4 5 OAI21D0BWP7T $T=217720 155000 1 180 $X=214630 $Y=154765
X832 230 227 192 34 4 5 OAI21D0BWP7T $T=226680 162840 1 180 $X=223590 $Y=162605
X833 50 229 32 221 4 5 OAI21D0BWP7T $T=245720 202040 1 180 $X=242630 $Y=201805
X834 272 274 246 276 4 5 OAI21D0BWP7T $T=273720 178520 1 0 $X=273430 $Y=174310
X835 309 315 314 34 4 5 OAI21D0BWP7T $T=316280 162840 0 180 $X=313190 $Y=158630
X836 290 332 257 328 4 5 OAI21D0BWP7T $T=334200 209880 0 0 $X=333910 $Y=209645
X837 67 345 277 340 4 5 OAI21D0BWP7T $T=340360 241240 1 0 $X=340070 $Y=237030
X838 80 81 83 84 4 5 OAI21D0BWP7T $T=352680 241240 1 0 $X=352390 $Y=237030
X839 85 363 86 378 4 5 OAI21D0BWP7T $T=357160 170680 1 0 $X=356870 $Y=166470
X840 85 361 87 359 4 5 OAI21D0BWP7T $T=360520 170680 1 180 $X=357430 $Y=170445
X841 85 369 96 368 4 5 OAI21D0BWP7T $T=374520 209880 0 0 $X=374230 $Y=209645
X842 85 375 97 372 4 5 OAI21D0BWP7T $T=377320 202040 0 0 $X=377030 $Y=201805
X843 85 374 98 377 4 5 OAI21D0BWP7T $T=377320 217720 1 0 $X=377030 $Y=213510
X844 85 376 101 365 4 5 OAI21D0BWP7T $T=381800 186360 0 180 $X=378710 $Y=182150
X845 99 100 102 103 4 5 OAI21D0BWP7T $T=379000 233400 0 0 $X=378710 $Y=233165
X846 97 383 104 381 4 5 OAI21D0BWP7T $T=390760 178520 1 180 $X=387670 $Y=178285
X847 96 384 104 387 4 5 OAI21D0BWP7T $T=392440 209880 0 0 $X=392150 $Y=209645
X848 87 393 104 390 4 5 OAI21D0BWP7T $T=393560 170680 1 0 $X=393270 $Y=166470
X849 106 385 99 388 4 5 OAI21D0BWP7T $T=398600 225560 1 180 $X=395510 $Y=225325
X850 85 382 108 389 4 5 OAI21D0BWP7T $T=399720 217720 0 0 $X=399430 $Y=217485
X851 101 394 104 401 4 5 OAI21D0BWP7T $T=408680 186360 1 0 $X=408390 $Y=182150
X852 98 396 104 399 4 5 OAI21D0BWP7T $T=408680 225560 1 0 $X=408390 $Y=221350
X853 83 392 102 110 4 5 OAI21D0BWP7T $T=408680 241240 1 0 $X=408390 $Y=237030
X854 85 397 109 398 4 5 OAI21D0BWP7T $T=412600 202040 0 180 $X=409510 $Y=197830
X855 86 406 104 395 4 5 OAI21D0BWP7T $T=418760 170680 1 180 $X=415670 $Y=170445
X856 109 407 104 409 4 5 OAI21D0BWP7T $T=417640 186360 1 0 $X=417350 $Y=182150
X857 108 410 104 403 4 5 OAI21D0BWP7T $T=421000 209880 0 180 $X=417910 $Y=205670
X858 116 411 86 412 4 5 OAI21D0BWP7T $T=423240 178520 0 0 $X=422950 $Y=178285
X859 116 414 87 419 4 5 OAI21D0BWP7T $T=432760 155000 0 0 $X=432470 $Y=154765
X860 116 413 101 416 4 5 OAI21D0BWP7T $T=434440 186360 1 0 $X=434150 $Y=182150
X861 116 415 96 421 4 5 OAI21D0BWP7T $T=436120 202040 0 0 $X=435830 $Y=201805
X862 116 122 109 417 4 5 OAI21D0BWP7T $T=441160 170680 1 180 $X=438070 $Y=170445
X863 116 418 108 125 4 5 OAI21D0BWP7T $T=441160 209880 1 0 $X=440870 $Y=205670
X864 116 420 98 124 4 5 OAI21D0BWP7T $T=444520 217720 1 180 $X=441430 $Y=217485
X895 17 4 10 20 5 149 ND3D0BWP7T $T=172360 162840 1 0 $X=172070 $Y=158630
X896 35 4 10 36 5 214 ND3D0BWP7T $T=214360 209880 1 0 $X=214070 $Y=205670
X897 246 4 52 61 5 276 ND3D0BWP7T $T=282680 186360 1 0 $X=282390 $Y=182150
X898 234 4 356 41 5 342 ND3D0BWP7T $T=360520 155000 1 180 $X=357430 $Y=154765
X899 4 5 DCAP16BWP7T $T=174040 209880 1 0 $X=173750 $Y=205670
X900 4 5 DCAP16BWP7T $T=180200 233400 1 0 $X=179910 $Y=229190
X901 4 5 DCAP16BWP7T $T=187480 155000 0 0 $X=187190 $Y=154765
X902 4 5 DCAP16BWP7T $T=198120 162840 0 0 $X=197830 $Y=162605
X903 4 5 DCAP16BWP7T $T=198120 170680 1 0 $X=197830 $Y=166470
X904 4 5 DCAP16BWP7T $T=206520 162840 1 0 $X=206230 $Y=158630
X905 4 5 DCAP16BWP7T $T=223320 178520 0 0 $X=223030 $Y=178285
X906 4 5 DCAP16BWP7T $T=229480 233400 1 0 $X=229190 $Y=229190
X907 4 5 DCAP16BWP7T $T=240120 186360 0 0 $X=239830 $Y=186125
X908 4 5 DCAP16BWP7T $T=240120 202040 1 0 $X=239830 $Y=197830
X909 4 5 DCAP16BWP7T $T=240120 241240 1 0 $X=239830 $Y=237030
X910 4 5 DCAP16BWP7T $T=251320 209880 0 0 $X=251030 $Y=209645
X911 4 5 DCAP16BWP7T $T=254680 225560 1 0 $X=254390 $Y=221350
X912 4 5 DCAP16BWP7T $T=271480 233400 0 0 $X=271190 $Y=233165
X913 4 5 DCAP16BWP7T $T=282120 178520 1 0 $X=281830 $Y=174310
X914 4 5 DCAP16BWP7T $T=282120 241240 1 0 $X=281830 $Y=237030
X915 4 5 DCAP16BWP7T $T=296120 170680 0 0 $X=295830 $Y=170445
X916 4 5 DCAP16BWP7T $T=324120 170680 0 0 $X=323830 $Y=170445
X917 4 5 DCAP16BWP7T $T=324120 209880 1 0 $X=323830 $Y=205670
X918 4 5 DCAP16BWP7T $T=324120 225560 0 0 $X=323830 $Y=225325
X919 4 5 DCAP16BWP7T $T=324120 233400 0 0 $X=323830 $Y=233165
X920 4 5 DCAP16BWP7T $T=324120 241240 1 0 $X=323830 $Y=237030
X921 4 5 DCAP16BWP7T $T=336440 217720 1 0 $X=336150 $Y=213510
X922 4 5 DCAP16BWP7T $T=342040 155000 0 0 $X=341750 $Y=154765
X923 4 5 DCAP16BWP7T $T=342040 170680 1 0 $X=341750 $Y=166470
X924 4 5 DCAP16BWP7T $T=343160 241240 1 0 $X=342870 $Y=237030
X925 4 5 DCAP16BWP7T $T=351000 202040 0 0 $X=350710 $Y=201805
X926 4 5 DCAP16BWP7T $T=355480 233400 1 0 $X=355190 $Y=229190
X927 4 5 DCAP16BWP7T $T=366120 155000 0 0 $X=365830 $Y=154765
X928 4 5 DCAP16BWP7T $T=366120 225560 1 0 $X=365830 $Y=221350
X929 4 5 DCAP16BWP7T $T=381800 178520 1 0 $X=381510 $Y=174310
X930 4 5 DCAP16BWP7T $T=381800 233400 0 0 $X=381510 $Y=233165
X931 4 5 DCAP16BWP7T $T=383480 225560 0 0 $X=383190 $Y=225325
X932 4 5 DCAP16BWP7T $T=384040 170680 1 0 $X=383750 $Y=166470
X933 4 5 DCAP16BWP7T $T=386840 194200 0 0 $X=386550 $Y=193965
X934 4 5 DCAP16BWP7T $T=389640 241240 1 0 $X=389350 $Y=237030
X935 4 5 DCAP16BWP7T $T=390760 178520 0 0 $X=390470 $Y=178285
X936 4 5 DCAP16BWP7T $T=390760 202040 1 0 $X=390470 $Y=197830
X937 4 5 DCAP16BWP7T $T=391320 233400 1 0 $X=391030 $Y=229190
X938 4 5 DCAP16BWP7T $T=392440 225560 1 0 $X=392150 $Y=221350
X939 4 5 DCAP16BWP7T $T=396360 155000 0 0 $X=396070 $Y=154765
X940 4 5 DCAP16BWP7T $T=398040 217720 1 0 $X=397750 $Y=213510
X941 4 5 DCAP16BWP7T $T=408120 209880 1 0 $X=407830 $Y=205670
X942 4 5 DCAP16BWP7T $T=420440 186360 1 0 $X=420150 $Y=182150
X943 4 5 DCAP16BWP7T $T=426040 202040 0 0 $X=425750 $Y=201805
X944 4 5 DCAP16BWP7T $T=432200 194200 0 0 $X=431910 $Y=193965
X970 22 4 134 19 168 5 NR3D1BWP7T $T=177960 202040 0 0 $X=177670 $Y=201805
X971 255 4 54 190 180 5 NR3D1BWP7T $T=253560 194200 1 0 $X=253270 $Y=189990
X972 255 4 62 208 250 5 NR3D1BWP7T $T=287160 202040 1 0 $X=286870 $Y=197830
X973 255 4 290 209 295 5 NR3D1BWP7T $T=296120 202040 1 0 $X=295830 $Y=197830
X974 174 171 4 5 172 173 MAOI222D1BWP7T $T=183000 194200 0 180 $X=178230 $Y=189990
X975 188 161 4 5 183 176 MAOI222D1BWP7T $T=190840 194200 0 180 $X=186070 $Y=189990
X976 314 303 4 5 310 325 MAOI222D1BWP7T $T=324680 162840 1 0 $X=324390 $Y=158630
X977 19 170 4 168 172 5 AOI21D1BWP7T $T=181880 202040 0 180 $X=178230 $Y=197830
X978 28 27 4 138 166 5 AOI21D1BWP7T $T=189160 217720 0 180 $X=185510 $Y=213510
X979 23 196 4 175 158 5 AOI21D1BWP7T $T=200360 217720 1 0 $X=200070 $Y=213510
X980 208 252 4 250 254 5 AOI21D1BWP7T $T=256360 194200 1 180 $X=252710 $Y=193965
X981 209 360 4 295 326 5 AOI21D1BWP7T $T=360520 178520 0 180 $X=356870 $Y=174310
X982 169 23 5 4 INVD2BWP7T $T=179640 162840 0 0 $X=179350 $Y=162605
X983 263 50 5 4 INVD2BWP7T $T=263640 225560 1 180 $X=261110 $Y=225325
X984 148 8 5 4 INVD2BWP7T $T=273160 225560 0 180 $X=270630 $Y=221350
X985 36 16 5 4 INVD2BWP7T $T=315720 225560 1 180 $X=313190 $Y=225325
X986 238 251 5 4 INVD2BWP7T $T=326920 202040 1 180 $X=324390 $Y=201805
X1020 24 177 4 5 169 DFQD0BWP7T $T=181880 162840 0 0 $X=181590 $Y=162605
X1021 24 215 4 5 200 DFQD0BWP7T $T=212120 170680 1 0 $X=211830 $Y=166470
X1022 24 222 4 5 17 DFQD0BWP7T $T=223320 178520 1 180 $X=212390 $Y=178285
X1023 24 236 4 5 197 DFQD0BWP7T $T=233960 186360 1 180 $X=223030 $Y=186125
X1024 24 213 4 5 157 DFQD0BWP7T $T=234520 162840 0 180 $X=223590 $Y=158630
X1025 24 229 4 5 35 DFQD0BWP7T $T=223880 202040 0 0 $X=223590 $Y=201805
X1026 24 245 4 5 249 DFQD0BWP7T $T=240680 162840 1 0 $X=240390 $Y=158630
X1027 24 244 4 5 246 DFQD0BWP7T $T=240680 178520 1 0 $X=240390 $Y=174310
X1028 24 243 4 5 195 DFQD0BWP7T $T=262520 170680 0 180 $X=251590 $Y=166470
X1029 24 258 4 5 247 DFQD0BWP7T $T=263080 209880 0 180 $X=252150 $Y=205670
X1030 24 268 4 5 212 DFQD0BWP7T $T=274840 162840 0 180 $X=263910 $Y=158630
X1031 24 201 4 5 189 DFQD0BWP7T $T=274840 225560 1 180 $X=263910 $Y=225325
X1032 24 63 4 5 278 DFQD0BWP7T $T=293320 233400 1 180 $X=282390 $Y=233165
X1033 24 64 4 5 263 DFQD0BWP7T $T=298360 225560 0 180 $X=287430 $Y=221350
X1034 24 296 4 5 307 DFQD0BWP7T $T=298920 162840 1 0 $X=298630 $Y=158630
X1035 69 308 4 5 299 DFQD0BWP7T $T=313480 225560 1 180 $X=302550 $Y=225325
X1036 69 374 4 5 89 DFQD0BWP7T $T=392440 225560 0 180 $X=381510 $Y=221350
X1037 69 383 4 5 373 DFQD0BWP7T $T=387960 186360 0 0 $X=387670 $Y=186125
X1038 69 392 4 5 105 DFQD0BWP7T $T=401960 233400 1 180 $X=391030 $Y=233165
X1039 69 393 4 5 371 DFQD0BWP7T $T=402520 162840 0 180 $X=391590 $Y=158630
X1040 69 394 4 5 366 DFQD0BWP7T $T=402520 178520 0 180 $X=391590 $Y=174310
X1041 69 384 4 5 370 DFQD0BWP7T $T=391880 202040 0 0 $X=391590 $Y=201805
X1042 69 406 4 5 380 DFQD0BWP7T $T=419320 162840 0 180 $X=408390 $Y=158630
X1043 69 396 4 5 379 DFQD0BWP7T $T=410360 225560 0 0 $X=410070 $Y=225325
X1044 69 386 4 5 111 DFQD0BWP7T $T=422680 241240 0 180 $X=411750 $Y=237030
X1045 69 397 4 5 356 DFQD0BWP7T $T=427160 202040 0 180 $X=416230 $Y=197830
X1046 69 410 4 5 391 DFQD0BWP7T $T=429400 209880 1 180 $X=418470 $Y=209645
X1047 69 411 4 5 400 DFQD0BWP7T $T=429960 162840 0 180 $X=419030 $Y=158630
X1048 69 407 4 5 408 DFQD0BWP7T $T=422680 170680 0 0 $X=422390 $Y=170445
X1049 69 413 4 5 404 DFQD0BWP7T $T=426040 186360 0 0 $X=425750 $Y=186125
X1050 69 415 4 5 402 DFQD0BWP7T $T=439480 202040 0 180 $X=428550 $Y=197830
X1051 69 414 4 5 405 DFQD0BWP7T $T=441160 162840 0 180 $X=430230 $Y=158630
X1052 69 418 4 5 112 DFQD0BWP7T $T=442280 217720 0 180 $X=431350 $Y=213510
X1053 69 420 4 5 113 DFQD0BWP7T $T=444520 225560 1 180 $X=433590 $Y=225325
X1054 69 123 4 5 118 DFQD0BWP7T $T=444520 241240 0 180 $X=433590 $Y=237030
X1055 25 26 4 5 INVD4BWP7T $T=183560 155000 0 0 $X=183270 $Y=154765
X1056 349 203 4 5 INVD4BWP7T $T=345400 233400 1 180 $X=341190 $Y=233165
X1057 23 4 5 8 22 178 NR3D0BWP7T $T=185800 209880 1 0 $X=185510 $Y=205670
X1058 27 4 5 14 22 141 NR3D0BWP7T $T=188600 241240 0 180 $X=185510 $Y=237030
X1059 256 4 5 251 255 288 NR3D0BWP7T $T=291080 162840 1 0 $X=290790 $Y=158630
X1060 180 5 192 190 194 4 AOI21D2BWP7T $T=187480 186360 0 0 $X=187190 $Y=186125
X1061 170 185 19 168 4 5 AOI21D0BWP7T $T=190840 202040 0 180 $X=187750 $Y=197830
X1062 230 243 192 227 4 5 AOI21D0BWP7T $T=243480 186360 0 180 $X=240390 $Y=182150
X1063 219 245 217 218 4 5 AOI21D0BWP7T $T=251880 155000 0 0 $X=251590 $Y=154765
X1064 235 275 256 271 4 5 AOI21D0BWP7T $T=275960 170680 1 180 $X=272870 $Y=170445
X1065 309 296 314 315 4 5 AOI21D0BWP7T $T=327480 162840 1 180 $X=324390 $Y=162605
X1066 178 4 5 175 BUFFD0BWP7T $T=188600 209880 1 0 $X=188310 $Y=205670
X1067 288 4 5 271 BUFFD0BWP7T $T=293880 162840 1 0 $X=293590 $Y=158630
X1068 385 4 5 386 BUFFD0BWP7T $T=393560 225560 0 0 $X=393270 $Y=225325
X1069 12 189 4 5 193 AN2D1BWP7T $T=189160 217720 1 0 $X=188870 $Y=213510
X1070 12 10 4 5 33 AN2D1BWP7T $T=216040 225560 1 180 $X=212950 $Y=225325
X1071 291 34 4 5 268 AN2D1BWP7T $T=298920 162840 0 180 $X=295830 $Y=158630
X1072 92 52 4 5 313 AN2D1BWP7T $T=369480 209880 0 180 $X=366390 $Y=205670
X1073 92 349 4 5 362 AN2D1BWP7T $T=369480 217720 1 180 $X=366390 $Y=217485
X1074 94 52 4 5 353 AN2D1BWP7T $T=373400 233400 0 180 $X=370310 $Y=229190
X1075 346 34 4 5 367 AN2D1BWP7T $T=375640 155000 0 0 $X=375350 $Y=154765
X1076 4 5 ICV_61 $T=198120 155000 0 0 $X=197830 $Y=154765
X1077 4 5 ICV_61 $T=198120 194200 1 0 $X=197830 $Y=189990
X1078 4 5 ICV_61 $T=198120 209880 1 0 $X=197830 $Y=205670
X1079 4 5 ICV_61 $T=198120 217720 0 0 $X=197830 $Y=217485
X1080 4 5 ICV_61 $T=198120 233400 0 0 $X=197830 $Y=233165
X1081 4 5 ICV_61 $T=226680 162840 0 0 $X=226390 $Y=162605
X1082 4 5 ICV_61 $T=226680 217720 1 0 $X=226390 $Y=213510
X1083 4 5 ICV_61 $T=240120 170680 1 0 $X=239830 $Y=166470
X1084 4 5 ICV_61 $T=240120 209880 1 0 $X=239830 $Y=205670
X1085 4 5 ICV_61 $T=262520 170680 1 0 $X=262230 $Y=166470
X1086 4 5 ICV_61 $T=324120 186360 1 0 $X=323830 $Y=182150
X1087 4 5 ICV_61 $T=366120 241240 1 0 $X=365830 $Y=237030
X1088 4 5 ICV_61 $T=380120 202040 0 0 $X=379830 $Y=201805
X1089 4 5 ICV_61 $T=395800 162840 0 0 $X=395510 $Y=162605
X1090 4 5 ICV_61 $T=422680 241240 1 0 $X=422390 $Y=237030
X1091 4 5 ICV_61 $T=426040 194200 1 0 $X=425750 $Y=189990
X1092 4 5 ICV_61 $T=428840 217720 0 0 $X=428550 $Y=217485
X1093 4 5 ICV_61 $T=437240 186360 1 0 $X=436950 $Y=182150
X1094 161 183 184 5 4 202 XOR3D0BWP7T $T=198680 178520 1 0 $X=198390 $Y=174310
X1095 174 185 171 5 4 204 XNR3D0BWP7T $T=199800 186360 0 0 $X=199510 $Y=186125
X1096 163 165 198 5 4 206 XNR3D0BWP7T $T=211000 194200 1 0 $X=210710 $Y=189990
X1097 32 209 4 206 5 215 31 OAI22D1BWP7T $T=211560 162840 1 180 $X=207350 $Y=162605
X1098 32 190 4 204 5 213 31 OAI22D1BWP7T $T=213240 178520 0 180 $X=209030 $Y=174310
X1099 163 198 4 216 199 5 IOA21D0BWP7T $T=211000 209880 1 0 $X=210710 $Y=205670
X1100 214 4 34 35 5 220 221 OAI211D0BWP7T $T=220520 209880 0 180 $X=216870 $Y=205670
X1101 234 34 231 39 4 5 226 AO22D0BWP7T $T=229480 178520 0 180 $X=224710 $Y=174310
X1102 44 239 192 233 4 5 MAOI222D2BWP7T $T=234520 209880 1 180 $X=226950 $Y=209645
X1103 217 260 259 266 4 5 MAOI222D2BWP7T $T=260280 170680 0 0 $X=259990 $Y=170445
X1104 24 226 4 5 47 DFQD1BWP7T $T=251320 209880 1 180 $X=240390 $Y=209645
X1105 24 58 4 5 262 DFQD1BWP7T $T=275400 217720 0 180 $X=264470 $Y=213510
X1106 69 367 4 5 234 DFQD1BWP7T $T=377880 162840 1 180 $X=366950 $Y=162605
X1107 69 361 4 5 355 DFQD1BWP7T $T=381800 178520 0 180 $X=370870 $Y=174310
X1108 69 376 4 5 238 DFQD1BWP7T $T=381800 186360 1 180 $X=370870 $Y=186125
X1109 69 369 4 5 95 DFQD1BWP7T $T=389640 241240 0 180 $X=378710 $Y=237030
X1110 69 363 4 5 364 DFQD1BWP7T $T=390200 162840 0 180 $X=379270 $Y=158630
X1111 69 375 4 5 280 DFQD1BWP7T $T=390760 202040 0 180 $X=379830 $Y=197830
X1112 69 382 4 5 349 DFQD1BWP7T $T=392440 209880 1 180 $X=381510 $Y=209645
X1113 34 162 4 5 32 236 208 MOAI22D0BWP7T $T=241800 194200 0 0 $X=241510 $Y=193965
X1114 39 246 4 5 181 222 31 MOAI22D0BWP7T $T=246840 194200 0 180 $X=242630 $Y=189990
X1115 48 144 240 248 53 4 5 XNR4D0BWP7T $T=241800 225560 1 0 $X=241510 $Y=221350
X1116 354 342 74 351 347 4 5 XNR4D0BWP7T $T=357720 186360 1 180 $X=344550 $Y=186125
X1117 358 82 352 341 337 4 5 XNR4D0BWP7T $T=358280 217720 0 180 $X=345110 $Y=213510
X1118 352 357 354 327 344 4 5 XNR4D0BWP7T $T=358840 202040 0 180 $X=345670 $Y=197830
X1119 247 148 4 5 BUFFD12BWP7T $T=245720 202040 0 0 $X=245430 $Y=201805
X1120 32 4 256 177 202 31 5 OAI22D2BWP7T $T=256920 186360 0 180 $X=249910 $Y=182150
X1121 57 56 248 241 225 4 5 XOR4D0BWP7T $T=267000 241240 0 180 $X=253830 $Y=237030
X1122 55 4 5 22 CKND1BWP7T $T=259160 225560 1 180 $X=257190 $Y=225325
X1123 44 239 230 44 4 239 5 IAO22D2BWP7T $T=264760 217720 0 180 $X=258310 $Y=213510
X1124 262 10 4 5 BUFFD1P5BWP7T $T=261960 209880 0 0 $X=261670 $Y=209645
X1125 355 52 4 5 BUFFD1P5BWP7T $T=351000 162840 1 0 $X=350710 $Y=158630
X1126 52 54 5 4 CKND2BWP7T $T=275960 241240 0 180 $X=273430 $Y=237030
X1127 251 5 9 258 4 NR2D0BWP7T $T=284920 202040 0 180 $X=282390 $Y=197830
X1128 273 259 5 260 4 264 219 AOI22D1BWP7T $T=288280 162840 0 180 $X=284070 $Y=158630
X1129 41 4 5 255 INVD3BWP7T $T=284920 186360 0 0 $X=284630 $Y=186125
X1130 278 4 5 66 CKBD1BWP7T $T=300600 233400 1 180 $X=298070 $Y=233165
X1131 299 4 5 40 CKBD1BWP7T $T=300600 225560 0 0 $X=300310 $Y=225325
X1132 68 281 4 5 INVD1P5BWP7T $T=307880 241240 1 0 $X=307590 $Y=237030
X1133 303 310 5 4 310 309 303 MAOI22D0BWP7T $T=313480 162840 0 180 $X=309270 $Y=158630
X1134 257 328 327 290 332 4 5 OAI31D1BWP7T $T=329160 202040 0 0 $X=328870 $Y=201805
X1135 277 340 344 67 345 4 5 OAI31D1BWP7T $T=339240 209880 0 0 $X=338950 $Y=209645
X1136 234 343 342 5 4 339 OA21D0BWP7T $T=342600 186360 0 180 $X=338950 $Y=182150
X1137 366 365 238 90 85 5 4 AOI22D0BWP7T $T=370040 186360 0 180 $X=366390 $Y=182150
X1138 370 368 95 90 85 5 4 AOI22D0BWP7T $T=376200 217720 1 180 $X=372550 $Y=217485
X1139 371 359 52 90 85 5 4 AOI22D0BWP7T $T=377320 170680 1 180 $X=373670 $Y=170445
X1140 373 372 280 90 85 5 4 AOI22D0BWP7T $T=377880 202040 0 180 $X=374230 $Y=197830
X1141 379 377 89 90 85 5 4 AOI22D0BWP7T $T=383480 225560 1 180 $X=379830 $Y=225325
X1142 380 378 364 90 85 5 4 AOI22D0BWP7T $T=387960 170680 1 180 $X=384310 $Y=170445
X1143 391 389 349 90 85 5 4 AOI22D0BWP7T $T=397480 217720 1 180 $X=393830 $Y=217485
X1144 104 381 90 373 107 5 4 AOI22D0BWP7T $T=396920 194200 0 0 $X=396630 $Y=193965
X1145 104 395 90 380 400 5 4 AOI22D0BWP7T $T=408680 170680 0 0 $X=408390 $Y=170445
X1146 104 387 90 370 402 5 4 AOI22D0BWP7T $T=408680 209880 0 0 $X=408390 $Y=209645
X1147 104 401 90 366 404 5 4 AOI22D0BWP7T $T=410920 186360 0 0 $X=410630 $Y=186125
X1148 408 398 356 90 85 5 4 AOI22D0BWP7T $T=414280 194200 1 180 $X=410630 $Y=193965
X1149 104 390 90 371 405 5 4 AOI22D0BWP7T $T=412600 178520 0 0 $X=412310 $Y=178285
X1150 104 403 90 391 112 5 4 AOI22D0BWP7T $T=412600 217720 1 0 $X=412310 $Y=213510
X1151 104 399 90 379 113 5 4 AOI22D0BWP7T $T=416520 217720 0 0 $X=416230 $Y=217485
X1152 104 409 90 408 115 5 4 AOI22D0BWP7T $T=419320 186360 0 0 $X=419030 $Y=186125
X1153 106 388 90 111 118 5 4 AOI22D0BWP7T $T=425480 217720 0 0 $X=425190 $Y=217485
X1154 106 117 90 119 120 5 4 AOI22D0BWP7T $T=426600 233400 1 0 $X=426310 $Y=229190
X1155 116 412 90 400 121 5 4 AOI22D0BWP7T $T=432200 178520 1 0 $X=431910 $Y=174310
X1156 116 416 90 404 128 5 4 AOI22D0BWP7T $T=438360 194200 1 0 $X=438070 $Y=189990
X1157 116 419 90 405 126 5 4 AOI22D0BWP7T $T=441160 162840 1 0 $X=440870 $Y=158630
X1158 116 417 90 115 129 5 4 AOI22D0BWP7T $T=441160 178520 1 0 $X=440870 $Y=174310
X1159 116 421 90 402 127 5 4 AOI22D0BWP7T $T=441160 202040 1 0 $X=440870 $Y=197830
X1160 114 5 69 4 CKND10BWP7T $T=422680 225560 0 0 $X=422390 $Y=225325
.ENDS
***************************************
.SUBCKT ICV_76 1 2
** N=2 EP=2 IP=4 FDC=24
*.SEEDPROM
X1 2 1 DCAP32BWP7T $T=1120 0 0 0 $X=830 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_41 1 2
** N=2 EP=2 IP=4 FDC=18
*.SEEDPROM
X0 1 2 DCAP8BWP7T $T=8960 0 0 0 $X=8670 $Y=-235
X1 1 2 DCAP16BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_37 1 2
** N=2 EP=2 IP=4 FDC=4
*.SEEDPROM
X0 1 2 DCAP4BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_60 1 2
** N=2 EP=2 IP=4 FDC=6
*.SEEDPROM
X1 1 2 DCAP8BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_43 1 2
** N=2 EP=2 IP=4 FDC=4
*.SEEDPROM
X1 1 2 DCAP4BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_55 1 2
** N=2 EP=2 IP=4 FDC=10
*.SEEDPROM
X0 1 2 ICV_40 $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_52 1 2
** N=2 EP=2 IP=4 FDC=6
*.SEEDPROM
X0 2 1 DCAPBWP7T $T=2240 0 0 0 $X=1950 $Y=-235
X1 1 2 DCAP4BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_54 1 2
** N=2 EP=2 IP=4 FDC=6
*.SEEDPROM
X0 1 2 DCAP8BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT NR2XD0BWP7T A2 VDD A1 ZN VSS
** N=6 EP=5 IP=0 FDC=4
*.SEEDPROM
M0 ZN A2 VSS VSS N L=1.8e-07 W=5e-07 $X=720 $Y=360 $D=0
M1 VSS A1 ZN VSS N L=1.8e-07 W=5e-07 $X=1440 $Y=360 $D=0
M2 6 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=720 $Y=2205 $D=16
M3 ZN A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=1320 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_38 1 2
** N=2 EP=2 IP=4 FDC=6
*.SEEDPROM
X1 1 2 DCAP8BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_45 1 2
** N=2 EP=2 IP=4 FDC=36
*.SEEDPROM
X0 2 1 DCAP32BWP7T $T=0 0 0 0 $X=-290 $Y=-235
X1 1 2 DCAP16BWP7T $T=17920 0 0 0 $X=17630 $Y=-235
.ENDS
***************************************
.SUBCKT INVD2P5BWP7T I ZN VSS VDD
** N=4 EP=4 IP=0 FDC=6
*.SEEDPROM
M0 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 VSS I ZN VSS N L=1.8e-07 W=4.65e-07 $X=2060 $Y=880 $D=0
M3 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M4 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M5 VDD I ZN VDD P L=1.8e-07 W=6.85e-07 $X=2060 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT BUFFD3BWP7T I VSS VDD Z
** N=5 EP=4 IP=0 FDC=8
*.SEEDPROM
M0 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=680 $Y=345 $D=0
M1 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=1570 $Y=345 $D=0
M2 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=2400 $Y=345 $D=0
M3 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=3120 $Y=345 $D=0
M4 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=680 $Y=2205 $D=16
M5 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1570 $Y=2205 $D=16
M6 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=2400 $Y=2205 $D=16
M7 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3120 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT BUFFD1BWP7T I VSS VDD Z
** N=5 EP=4 IP=0 FDC=4
*.SEEDPROM
M0 VSS I 5 VSS N L=1.8e-07 W=5e-07 $X=625 $Y=845 $D=0
M1 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=1425 $Y=345 $D=0
M2 VDD I 5 VDD P L=1.8e-07 W=6.85e-07 $X=625 $Y=2205 $D=16
M3 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1425 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IAO21D0BWP7T A1 A2 VSS VDD B ZN
** N=9 EP=6 IP=0 FDC=8
*.SEEDPROM
M0 7 A1 VSS VSS N L=1.8e-07 W=4.2e-07 $X=460 $Y=730 $D=0
M1 VSS A2 7 VSS N L=1.8e-07 W=4.2e-07 $X=1180 $Y=730 $D=0
M2 ZN 7 VSS VSS N L=1.8e-07 W=5e-07 $X=1900 $Y=730 $D=0
M3 VSS B ZN VSS N L=1.8e-07 W=5e-07 $X=2620 $Y=730 $D=0
M4 8 A1 7 VDD P L=1.8e-07 W=4.2e-07 $X=620 $Y=2860 $D=16
M5 VDD A2 8 VDD P L=1.8e-07 W=4.2e-07 $X=1185 $Y=2860 $D=16
M6 9 7 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1945 $Y=2860 $D=16
M7 ZN B 9 VDD P L=1.8e-07 W=6.85e-07 $X=2515 $Y=2860 $D=16
.ENDS
***************************************
.SUBCKT AN3D1BWP7T A1 A2 A3 VDD VSS Z
** N=9 EP=6 IP=0 FDC=8
*.SEEDPROM
M0 8 A1 7 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=345 $D=0
M1 9 A2 8 VSS N L=1.8e-07 W=5e-07 $X=1205 $Y=345 $D=0
M2 VSS A3 9 VSS N L=1.8e-07 W=5e-07 $X=1790 $Y=345 $D=0
M3 Z 7 VSS VSS N L=1.8e-07 W=1e-06 $X=2560 $Y=345 $D=0
M4 VDD A1 7 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2205 $D=16
M5 7 A2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1230 $Y=2205 $D=16
M6 VDD A3 7 VDD P L=1.8e-07 W=6.85e-07 $X=1950 $Y=2205 $D=16
M7 Z 7 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2560 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INVD12BWP7T I ZN VSS VDD
** N=4 EP=4 IP=0 FDC=24
*.SEEDPROM
M0 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=2060 $Y=345 $D=0
M3 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=2780 $Y=345 $D=0
M4 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=3520 $Y=345 $D=0
M5 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=4240 $Y=345 $D=0
M6 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=4970 $Y=345 $D=0
M7 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=5690 $Y=345 $D=0
M8 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=6450 $Y=345 $D=0
M9 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=7170 $Y=345 $D=0
M10 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=7890 $Y=345 $D=0
M11 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=8650 $Y=345 $D=0
M12 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M13 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M14 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M15 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M16 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=3520 $Y=2205 $D=16
M17 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=4240 $Y=2205 $D=16
M18 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=4970 $Y=2205 $D=16
M19 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=5690 $Y=2205 $D=16
M20 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=6450 $Y=2205 $D=16
M21 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=7170 $Y=2205 $D=16
M22 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=7890 $Y=2205 $D=16
M23 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=8650 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKND12BWP7T I VDD ZN VSS
** N=4 EP=4 IP=0 FDC=22
*.SEEDPROM
M0 ZN I VSS VSS N L=1.8e-07 W=6.3e-07 $X=1340 $Y=410 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=6.3e-07 $X=2060 $Y=410 $D=0
M2 ZN I VSS VSS N L=1.8e-07 W=6.3e-07 $X=2780 $Y=410 $D=0
M3 VSS I ZN VSS N L=1.8e-07 W=6.3e-07 $X=3500 $Y=410 $D=0
M4 ZN I VSS VSS N L=1.8e-07 W=6.3e-07 $X=4220 $Y=410 $D=0
M5 VSS I ZN VSS N L=1.8e-07 W=6.3e-07 $X=4940 $Y=410 $D=0
M6 ZN I VSS VSS N L=1.8e-07 W=6.3e-07 $X=5660 $Y=410 $D=0
M7 VSS I ZN VSS N L=1.8e-07 W=6.3e-07 $X=6380 $Y=410 $D=0
M8 ZN I VSS VSS N L=1.8e-07 W=6.3e-07 $X=7100 $Y=410 $D=0
M9 VSS I ZN VSS N L=1.8e-07 W=6.3e-07 $X=7820 $Y=410 $D=0
M10 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M11 VDD I ZN VDD P L=1.8e-07 W=1.525e-06 $X=1340 $Y=2050 $D=16
M12 ZN I VDD VDD P L=1.8e-07 W=1.525e-06 $X=2060 $Y=2050 $D=16
M13 VDD I ZN VDD P L=1.8e-07 W=1.525e-06 $X=2780 $Y=2050 $D=16
M14 ZN I VDD VDD P L=1.8e-07 W=1.525e-06 $X=3500 $Y=2050 $D=16
M15 VDD I ZN VDD P L=1.8e-07 W=1.525e-06 $X=4220 $Y=2050 $D=16
M16 ZN I VDD VDD P L=1.8e-07 W=1.525e-06 $X=4940 $Y=2050 $D=16
M17 VDD I ZN VDD P L=1.8e-07 W=1.525e-06 $X=5660 $Y=2050 $D=16
M18 ZN I VDD VDD P L=1.8e-07 W=1.525e-06 $X=6380 $Y=2050 $D=16
M19 VDD I ZN VDD P L=1.8e-07 W=1.525e-06 $X=7100 $Y=2050 $D=16
M20 ZN I VDD VDD P L=1.8e-07 W=1.345e-06 $X=7820 $Y=2230 $D=16
D21 VSS I DN AREA=2.037e-13 PJ=1.81e-06 $X=140 $Y=645 $D=32
.ENDS
***************************************
.SUBCKT DFQD2BWP7T CP D Q VSS VDD
** N=16 EP=5 IP=0 FDC=26
*.SEEDPROM
M0 VSS CP 6 VSS N L=1.8e-07 W=5e-07 $X=640 $Y=840 $D=0
M1 9 6 VSS VSS N L=1.8e-07 W=5e-07 $X=1240 $Y=840 $D=0
M2 13 6 VSS VSS N L=1.8e-07 W=9.4e-07 $X=2665 $Y=405 $D=0
M3 7 D 13 VSS N L=1.8e-07 W=9.4e-07 $X=3135 $Y=405 $D=0
M4 14 9 7 VSS N L=1.8e-07 W=4.2e-07 $X=3990 $Y=895 $D=0
M5 VSS 8 14 VSS N L=1.8e-07 W=4.2e-07 $X=4485 $Y=895 $D=0
M6 8 7 VSS VSS N L=1.8e-07 W=5.4e-07 $X=5285 $Y=775 $D=0
M7 11 9 8 VSS N L=1.8e-07 W=9.1e-07 $X=6005 $Y=405 $D=0
M8 10 6 11 VSS N L=1.8e-07 W=4.2e-07 $X=6725 $Y=895 $D=0
M9 VSS 12 10 VSS N L=1.8e-07 W=4.2e-07 $X=7445 $Y=895 $D=0
M10 12 11 VSS VSS N L=1.8e-07 W=1e-06 $X=8235 $Y=345 $D=0
M11 Q 12 VSS VSS N L=1.8e-07 W=1e-06 $X=9680 $Y=345 $D=0
M12 VSS 12 Q VSS N L=1.8e-07 W=1e-06 $X=10400 $Y=345 $D=0
M13 VDD CP 6 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2345 $D=16
M14 9 6 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1240 $Y=2345 $D=16
M15 15 9 VDD VDD P L=1.8e-07 W=9.2e-07 $X=2705 $Y=2205 $D=16
M16 7 D 15 VDD P L=1.8e-07 W=9.2e-07 $X=3205 $Y=2205 $D=16
M17 16 6 7 VDD P L=1.8e-07 W=4.2e-07 $X=3985 $Y=2705 $D=16
M18 VDD 8 16 VDD P L=1.8e-07 W=4.2e-07 $X=4485 $Y=2705 $D=16
M19 8 7 VDD VDD P L=1.8e-07 W=9.6e-07 $X=5285 $Y=2175 $D=16
M20 11 6 8 VDD P L=1.8e-07 W=1.34e-06 $X=6005 $Y=2175 $D=16
M21 10 9 11 VDD P L=1.8e-07 W=4.2e-07 $X=6725 $Y=2470 $D=16
M22 VDD 12 10 VDD P L=1.8e-07 W=4.2e-07 $X=7485 $Y=2205 $D=16
M23 12 11 VDD VDD P L=1.8e-07 W=1.37e-06 $X=8260 $Y=2205 $D=16
M24 Q 12 VDD VDD P L=1.8e-07 W=1.37e-06 $X=9680 $Y=2205 $D=16
M25 VDD 12 Q VDD P L=1.8e-07 W=1.37e-06 $X=10400 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT BUFFD5BWP7T I VSS VDD Z
** N=5 EP=4 IP=0 FDC=14
*.SEEDPROM
M0 5 I VSS VSS N L=1.8e-07 W=1e-06 $X=640 $Y=345 $D=0
M1 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=1360 $Y=345 $D=0
M2 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=2140 $Y=345 $D=0
M3 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=2860 $Y=345 $D=0
M4 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=3640 $Y=345 $D=0
M5 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=4360 $Y=345 $D=0
M6 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=5140 $Y=345 $D=0
M7 5 I VDD VDD P L=1.8e-07 W=1.37e-06 $X=640 $Y=2205 $D=16
M8 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=1360 $Y=2205 $D=16
M9 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2140 $Y=2205 $D=16
M10 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=2860 $Y=2205 $D=16
M11 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3640 $Y=2205 $D=16
M12 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=4360 $Y=2205 $D=16
M13 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=5140 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT BUFFD2BWP7T I Z VSS VDD
** N=5 EP=4 IP=0 FDC=6
*.SEEDPROM
M0 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=680 $Y=345 $D=0
M1 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=1590 $Y=345 $D=0
M2 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=2430 $Y=345 $D=0
M3 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=680 $Y=2205 $D=16
M4 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1590 $Y=2205 $D=16
M5 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=2430 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ND2D2BWP7T A1 ZN A2 VSS VDD
** N=7 EP=5 IP=0 FDC=8
*.SEEDPROM
M0 6 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=700 $Y=345 $D=0
M1 ZN A1 6 VSS N L=1.8e-07 W=1e-06 $X=1420 $Y=345 $D=0
M2 7 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=2260 $Y=345 $D=0
M3 VSS A2 7 VSS N L=1.8e-07 W=1e-06 $X=2980 $Y=345 $D=0
M4 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=700 $Y=2205 $D=16
M5 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1420 $Y=2205 $D=16
M6 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2260 $Y=2205 $D=16
M7 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2980 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKND2D2BWP7T A2 VSS A1 ZN VDD
** N=6 EP=5 IP=0 FDC=8
*.SEEDPROM
M0 VSS A2 6 VSS N L=1.8e-07 W=6e-07 $X=660 $Y=545 $D=0
M1 6 A2 VSS VSS N L=1.8e-07 W=6e-07 $X=1380 $Y=545 $D=0
M2 ZN A1 6 VSS N L=1.8e-07 W=8e-07 $X=2320 $Y=545 $D=0
M3 6 A1 ZN VSS N L=1.8e-07 W=8e-07 $X=3120 $Y=545 $D=0
M4 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M5 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1380 $Y=2205 $D=16
M6 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2320 $Y=2205 $D=16
M7 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3120 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ND2D1P5BWP7T A1 ZN A2 VSS VDD
** N=7 EP=5 IP=0 FDC=8
*.SEEDPROM
M0 6 A2 VSS VSS N L=1.8e-07 W=7.5e-07 $X=740 $Y=345 $D=0
M1 ZN A1 6 VSS N L=1.8e-07 W=7.5e-07 $X=1360 $Y=345 $D=0
M2 7 A1 ZN VSS N L=1.8e-07 W=7.5e-07 $X=2080 $Y=345 $D=0
M3 VSS A2 7 VSS N L=1.8e-07 W=7.5e-07 $X=2690 $Y=345 $D=0
M4 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=740 $Y=2205 $D=16
M5 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1460 $Y=2205 $D=16
M6 ZN A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=2260 $Y=2205 $D=16
M7 VDD A2 ZN VDD P L=1.8e-07 W=6.85e-07 $X=2980 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_83 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244
** N=595 EP=242 IP=4232 FDC=11015
*.SEEDPROM
M0 37 46 3 3 N L=1.8e-07 W=1e-06 $X=204360 $Y=257265 $D=0
M1 3 46 37 3 N L=1.8e-07 W=1e-06 $X=205080 $Y=257265 $D=0
M2 37 46 3 3 N L=1.8e-07 W=1e-06 $X=205800 $Y=257265 $D=0
M3 3 46 37 3 N L=1.8e-07 W=1e-06 $X=206520 $Y=257265 $D=0
M4 37 46 3 3 N L=1.8e-07 W=1e-06 $X=207240 $Y=257265 $D=0
M5 3 46 37 3 N L=1.8e-07 W=1e-06 $X=207960 $Y=257265 $D=0
M6 69 11 3 3 N L=1.8e-07 W=7e-07 $X=296920 $Y=280785 $D=0
M7 3 11 69 3 N L=1.8e-07 W=7e-07 $X=297720 $Y=280785 $D=0
M8 69 11 3 3 N L=1.8e-07 W=7e-07 $X=298440 $Y=280785 $D=0
M9 595 147 145 3 N L=1.8e-07 W=1e-06 $X=330025 $Y=257265 $D=0
M10 3 472 595 3 N L=1.8e-07 W=1e-06 $X=330760 $Y=257265 $D=0
M11 145 151 3 3 N L=1.8e-07 W=1e-06 $X=331720 $Y=257265 $D=0
M12 3 35 145 3 N L=1.8e-07 W=1e-06 $X=332850 $Y=257265 $D=0
M13 37 46 4 4 P L=1.8e-07 W=1.37e-06 $X=204360 $Y=259125 $D=16
M14 4 46 37 4 P L=1.8e-07 W=1.37e-06 $X=205080 $Y=259125 $D=16
M15 37 46 4 4 P L=1.8e-07 W=1.37e-06 $X=205800 $Y=259125 $D=16
M16 4 46 37 4 P L=1.8e-07 W=1.37e-06 $X=206520 $Y=259125 $D=16
M17 37 46 4 4 P L=1.8e-07 W=1.37e-06 $X=207240 $Y=259125 $D=16
M18 4 46 37 4 P L=1.8e-07 W=1.37e-06 $X=207960 $Y=259125 $D=16
M19 69 11 4 4 P L=1.8e-07 W=1.37e-06 $X=296920 $Y=282645 $D=16
M20 4 11 69 4 P L=1.8e-07 W=1.37e-06 $X=297640 $Y=282645 $D=16
M21 69 11 4 4 P L=1.8e-07 W=1.37e-06 $X=298440 $Y=282645 $D=16
M22 4 11 69 4 P L=1.8e-07 W=1.37e-06 $X=299160 $Y=282645 $D=16
M23 145 472 478 4 P L=1.8e-07 W=1.37e-06 $X=328695 $Y=259125 $D=16
M24 478 147 145 4 P L=1.8e-07 W=1.37e-06 $X=329420 $Y=259125 $D=16
M25 145 147 478 4 P L=1.8e-07 W=1.37e-06 $X=330220 $Y=259125 $D=16
M26 478 472 145 4 P L=1.8e-07 W=1.37e-06 $X=331000 $Y=259125 $D=16
M27 479 151 478 4 P L=1.8e-07 W=1.37e-06 $X=331720 $Y=259125 $D=16
M28 4 35 479 4 P L=1.8e-07 W=1.37e-06 $X=332440 $Y=259125 $D=16
M29 479 35 4 4 P L=1.8e-07 W=1.37e-06 $X=333240 $Y=259125 $D=16
M30 478 151 479 4 P L=1.8e-07 W=1.37e-06 $X=333960 $Y=259125 $D=16
D31 3 11 DN AREA=2.037e-13 PJ=1.81e-06 $X=299480 $Y=281300 $D=32
X223 4 3 DCAPBWP7T $T=162840 327480 1 0 $X=162550 $Y=323270
X224 4 3 DCAPBWP7T $T=162840 343160 1 0 $X=162550 $Y=338950
X225 4 3 DCAPBWP7T $T=167320 343160 0 0 $X=167030 $Y=342925
X226 4 3 DCAPBWP7T $T=171800 358840 1 0 $X=171510 $Y=354630
X227 4 3 DCAPBWP7T $T=173480 272600 1 0 $X=173190 $Y=268390
X228 4 3 DCAPBWP7T $T=177960 319640 1 0 $X=177670 $Y=315430
X229 4 3 DCAPBWP7T $T=195320 249080 1 0 $X=195030 $Y=244870
X230 4 3 DCAPBWP7T $T=195320 249080 0 0 $X=195030 $Y=248845
X231 4 3 DCAPBWP7T $T=195320 256920 1 0 $X=195030 $Y=252710
X232 4 3 DCAPBWP7T $T=195320 264760 0 0 $X=195030 $Y=264525
X233 4 3 DCAPBWP7T $T=198120 311800 1 0 $X=197830 $Y=307590
X234 4 3 DCAPBWP7T $T=213800 327480 1 0 $X=213510 $Y=323270
X235 4 3 DCAPBWP7T $T=219400 264760 1 0 $X=219110 $Y=260550
X236 4 3 DCAPBWP7T $T=237320 264760 1 0 $X=237030 $Y=260550
X237 4 3 DCAPBWP7T $T=237320 264760 0 0 $X=237030 $Y=264525
X238 4 3 DCAPBWP7T $T=237320 272600 1 0 $X=237030 $Y=268390
X239 4 3 DCAPBWP7T $T=237320 351000 0 0 $X=237030 $Y=350765
X240 4 3 DCAPBWP7T $T=240120 272600 1 0 $X=239830 $Y=268390
X241 4 3 DCAPBWP7T $T=251320 288280 1 0 $X=251030 $Y=284070
X242 4 3 DCAPBWP7T $T=253560 319640 0 0 $X=253270 $Y=319405
X243 4 3 DCAPBWP7T $T=253560 358840 1 0 $X=253270 $Y=354630
X244 4 3 DCAPBWP7T $T=264760 327480 0 0 $X=264470 $Y=327245
X245 4 3 DCAPBWP7T $T=267000 311800 0 0 $X=266710 $Y=311565
X246 4 3 DCAPBWP7T $T=272040 296120 0 0 $X=271750 $Y=295885
X247 4 3 DCAPBWP7T $T=291080 241240 0 0 $X=290790 $Y=241005
X248 4 3 DCAPBWP7T $T=302840 335320 0 0 $X=302550 $Y=335085
X249 4 3 DCAPBWP7T $T=307880 335320 0 0 $X=307590 $Y=335085
X250 4 3 DCAPBWP7T $T=310120 335320 1 0 $X=309830 $Y=331110
X251 4 3 DCAPBWP7T $T=321320 256920 1 0 $X=321030 $Y=252710
X252 4 3 DCAPBWP7T $T=321320 280440 1 0 $X=321030 $Y=276230
X253 4 3 DCAPBWP7T $T=321320 327480 1 0 $X=321030 $Y=323270
X254 4 3 DCAPBWP7T $T=321320 343160 0 0 $X=321030 $Y=342925
X255 4 3 DCAPBWP7T $T=328040 303960 0 0 $X=327750 $Y=303725
X256 4 3 DCAPBWP7T $T=338120 264760 0 0 $X=337830 $Y=264525
X257 4 3 DCAPBWP7T $T=355480 311800 0 0 $X=355190 $Y=311565
X258 4 3 DCAPBWP7T $T=363320 351000 1 0 $X=363030 $Y=346790
X259 4 3 DCAPBWP7T $T=366120 335320 1 0 $X=365830 $Y=331110
X260 4 3 DCAPBWP7T $T=384040 327480 1 0 $X=383750 $Y=323270
X261 4 3 DCAPBWP7T $T=387960 272600 0 0 $X=387670 $Y=272365
X262 4 3 DCAPBWP7T $T=397480 288280 1 0 $X=397190 $Y=284070
X263 4 3 DCAPBWP7T $T=405320 288280 0 0 $X=405030 $Y=288045
X264 4 3 DCAPBWP7T $T=405320 319640 1 0 $X=405030 $Y=315430
X265 4 3 DCAPBWP7T $T=405320 319640 0 0 $X=405030 $Y=319405
X266 4 3 DCAPBWP7T $T=405320 327480 0 0 $X=405030 $Y=327245
X267 4 3 DCAPBWP7T $T=405320 351000 0 0 $X=405030 $Y=350765
X268 4 3 DCAPBWP7T $T=408120 272600 0 0 $X=407830 $Y=272365
X269 4 3 DCAPBWP7T $T=408120 296120 1 0 $X=407830 $Y=291910
X270 4 3 DCAPBWP7T $T=408120 327480 1 0 $X=407830 $Y=323270
X271 4 3 DCAPBWP7T $T=414840 303960 0 0 $X=414550 $Y=303725
X272 4 3 DCAPBWP7T $T=421560 351000 1 0 $X=421270 $Y=346790
X273 4 3 DCAPBWP7T $T=430520 343160 0 0 $X=430230 $Y=342925
X274 4 3 DCAPBWP7T $T=430520 358840 1 0 $X=430230 $Y=354630
X275 4 3 DCAPBWP7T $T=435560 327480 0 0 $X=435270 $Y=327245
X276 4 3 DCAPBWP7T $T=437800 311800 0 0 $X=437510 $Y=311565
X277 4 3 DCAPBWP7T $T=447320 303960 0 0 $X=447030 $Y=303725
X278 4 3 DCAPBWP7T $T=447320 327480 1 0 $X=447030 $Y=323270
X279 4 3 DCAPBWP7T $T=447320 343160 0 0 $X=447030 $Y=342925
X280 4 3 DCAPBWP7T $T=447320 358840 1 0 $X=447030 $Y=354630
X281 3 4 DCAP8BWP7T $T=156120 351000 0 0 $X=155830 $Y=350765
X282 3 4 DCAP8BWP7T $T=158360 327480 1 0 $X=158070 $Y=323270
X283 3 4 DCAP8BWP7T $T=191960 319640 0 0 $X=191670 $Y=319405
X284 3 4 DCAP8BWP7T $T=192520 343160 1 0 $X=192230 $Y=338950
X285 3 4 DCAP8BWP7T $T=198120 264760 0 0 $X=197830 $Y=264525
X286 3 4 DCAP8BWP7T $T=225560 249080 0 0 $X=225270 $Y=248845
X287 3 4 DCAP8BWP7T $T=232840 272600 1 0 $X=232550 $Y=268390
X288 3 4 DCAP8BWP7T $T=233960 272600 0 0 $X=233670 $Y=272365
X289 3 4 DCAP8BWP7T $T=234520 335320 0 0 $X=234230 $Y=335085
X290 3 4 DCAP8BWP7T $T=234520 351000 1 0 $X=234230 $Y=346790
X291 3 4 DCAP8BWP7T $T=275960 319640 0 0 $X=275670 $Y=319405
X292 3 4 DCAP8BWP7T $T=276520 264760 0 0 $X=276230 $Y=264525
X293 3 4 DCAP8BWP7T $T=276520 327480 1 0 $X=276230 $Y=323270
X294 3 4 DCAP8BWP7T $T=317960 319640 1 0 $X=317670 $Y=315430
X295 3 4 DCAP8BWP7T $T=317960 351000 1 0 $X=317670 $Y=346790
X296 3 4 DCAP8BWP7T $T=318520 296120 1 0 $X=318230 $Y=291910
X297 3 4 DCAP8BWP7T $T=318520 311800 1 0 $X=318230 $Y=307590
X298 3 4 DCAP8BWP7T $T=318520 319640 0 0 $X=318230 $Y=319405
X299 3 4 DCAP8BWP7T $T=324120 335320 1 0 $X=323830 $Y=331110
X300 3 4 DCAP8BWP7T $T=340920 327480 0 0 $X=340630 $Y=327245
X301 3 4 DCAP8BWP7T $T=359960 241240 0 0 $X=359670 $Y=241005
X302 3 4 DCAP8BWP7T $T=360520 249080 1 0 $X=360230 $Y=244870
X303 3 4 DCAP8BWP7T $T=360520 343160 0 0 $X=360230 $Y=342925
X304 3 4 DCAP8BWP7T $T=366120 358840 1 0 $X=365830 $Y=354630
X305 3 4 DCAP8BWP7T $T=402520 288280 1 0 $X=402230 $Y=284070
X306 3 4 DCAP8BWP7T $T=402520 343160 0 0 $X=402230 $Y=342925
X307 3 4 DCAP8BWP7T $T=402520 351000 1 0 $X=402230 $Y=346790
X308 3 4 DCAP8BWP7T $T=426040 343160 0 0 $X=425750 $Y=342925
X309 3 4 DCAP8BWP7T $T=426040 358840 1 0 $X=425750 $Y=354630
X310 3 4 DCAP8BWP7T $T=431080 327480 0 0 $X=430790 $Y=327245
X311 3 4 DCAP8BWP7T $T=442840 358840 1 0 $X=442550 $Y=354630
X312 3 4 DCAP8BWP7T $T=444520 249080 0 0 $X=444230 $Y=248845
X313 3 4 DCAP8BWP7T $T=444520 256920 1 0 $X=444230 $Y=252710
X314 3 4 DCAP8BWP7T $T=444520 280440 1 0 $X=444230 $Y=276230
X315 3 4 DCAP8BWP7T $T=444520 288280 0 0 $X=444230 $Y=288045
X316 3 4 DCAP8BWP7T $T=444520 335320 0 0 $X=444230 $Y=335085
X317 3 4 DCAP4BWP7T $T=156120 288280 1 0 $X=155830 $Y=284070
X318 3 4 DCAP4BWP7T $T=172920 241240 0 0 $X=172630 $Y=241005
X319 3 4 DCAP4BWP7T $T=194200 351000 1 0 $X=193910 $Y=346790
X320 3 4 DCAP4BWP7T $T=194760 272600 1 0 $X=194470 $Y=268390
X321 3 4 DCAP4BWP7T $T=194760 311800 1 0 $X=194470 $Y=307590
X322 3 4 DCAP4BWP7T $T=236200 319640 0 0 $X=235910 $Y=319405
X323 3 4 DCAP4BWP7T $T=236760 296120 1 0 $X=236470 $Y=291910
X324 3 4 DCAP4BWP7T $T=240120 296120 1 0 $X=239830 $Y=291910
X325 3 4 DCAP4BWP7T $T=240120 303960 0 0 $X=239830 $Y=303725
X326 3 4 DCAP4BWP7T $T=249080 311800 1 0 $X=248790 $Y=307590
X327 3 4 DCAP4BWP7T $T=262520 335320 0 0 $X=262230 $Y=335085
X328 3 4 DCAP4BWP7T $T=266440 343160 1 0 $X=266150 $Y=338950
X329 3 4 DCAP4BWP7T $T=278200 256920 1 0 $X=277910 $Y=252710
X330 3 4 DCAP4BWP7T $T=278200 319640 1 0 $X=277910 $Y=315430
X331 3 4 DCAP4BWP7T $T=278200 358840 1 0 $X=277910 $Y=354630
X332 3 4 DCAP4BWP7T $T=278760 303960 0 0 $X=278470 $Y=303725
X333 3 4 DCAP4BWP7T $T=291080 296120 0 0 $X=290790 $Y=295885
X334 3 4 DCAP4BWP7T $T=291080 303960 0 0 $X=290790 $Y=303725
X335 3 4 DCAP4BWP7T $T=292760 264760 1 0 $X=292470 $Y=260550
X336 3 4 DCAP4BWP7T $T=320200 288280 1 0 $X=319910 $Y=284070
X337 3 4 DCAP4BWP7T $T=320760 249080 0 0 $X=320470 $Y=248845
X338 3 4 DCAP4BWP7T $T=320760 335320 0 0 $X=320470 $Y=335085
X339 3 4 DCAP4BWP7T $T=347080 264760 0 0 $X=346790 $Y=264525
X340 3 4 DCAP4BWP7T $T=384040 288280 1 0 $X=383750 $Y=284070
X341 3 4 DCAP4BWP7T $T=384040 296120 1 0 $X=383750 $Y=291910
X342 3 4 DCAP4BWP7T $T=395240 319640 1 0 $X=394950 $Y=315430
X343 3 4 DCAP4BWP7T $T=404200 241240 0 0 $X=403910 $Y=241005
X344 3 4 DCAP4BWP7T $T=404760 272600 0 0 $X=404470 $Y=272365
X345 3 4 DCAP4BWP7T $T=408120 319640 1 0 $X=407830 $Y=315430
X346 3 4 DCAP4BWP7T $T=429960 249080 0 0 $X=429670 $Y=248845
X347 3 4 DCAP4BWP7T $T=446760 280440 0 0 $X=446470 $Y=280205
X348 3 4 ICV_40 $T=156120 343160 1 0 $X=155830 $Y=338950
X349 3 4 ICV_40 $T=166760 272600 1 0 $X=166470 $Y=268390
X350 3 4 ICV_40 $T=169560 296120 0 0 $X=169270 $Y=295885
X351 3 4 ICV_40 $T=175720 288280 1 0 $X=175430 $Y=284070
X352 3 4 ICV_40 $T=190280 280440 0 0 $X=189990 $Y=280205
X353 3 4 ICV_40 $T=190280 296120 0 0 $X=189990 $Y=295885
X354 3 4 ICV_40 $T=190280 303960 0 0 $X=189990 $Y=303725
X355 3 4 ICV_40 $T=207080 327480 1 0 $X=206790 $Y=323270
X356 3 4 ICV_40 $T=231720 280440 1 0 $X=231430 $Y=276230
X357 3 4 ICV_40 $T=231720 280440 0 0 $X=231430 $Y=280205
X358 3 4 ICV_40 $T=249080 327480 1 0 $X=248790 $Y=323270
X359 3 4 ICV_40 $T=258040 303960 1 0 $X=257750 $Y=299750
X360 3 4 ICV_40 $T=258040 327480 0 0 $X=257750 $Y=327245
X361 3 4 ICV_40 $T=273720 272600 1 0 $X=273430 $Y=268390
X362 3 4 ICV_40 $T=273720 280440 0 0 $X=273430 $Y=280205
X363 3 4 ICV_40 $T=273720 296120 1 0 $X=273430 $Y=291910
X364 3 4 ICV_40 $T=282120 264760 1 0 $X=281830 $Y=260550
X365 3 4 ICV_40 $T=291080 272600 1 0 $X=290790 $Y=268390
X366 3 4 ICV_40 $T=298920 256920 0 0 $X=298630 $Y=256685
X367 3 4 ICV_40 $T=314600 280440 1 0 $X=314310 $Y=276230
X368 3 4 ICV_40 $T=315720 351000 0 0 $X=315430 $Y=350765
X369 3 4 ICV_40 $T=324120 343160 1 0 $X=323830 $Y=338950
X370 3 4 ICV_40 $T=342040 319640 1 0 $X=341750 $Y=315430
X371 3 4 ICV_40 $T=346520 256920 0 0 $X=346230 $Y=256685
X372 3 4 ICV_40 $T=350440 288280 0 0 $X=350150 $Y=288045
X373 3 4 ICV_40 $T=357720 319640 1 0 $X=357430 $Y=315430
X374 3 4 ICV_40 $T=358280 256920 1 0 $X=357990 $Y=252710
X375 3 4 ICV_40 $T=358280 256920 0 0 $X=357990 $Y=256685
X376 3 4 ICV_40 $T=358280 280440 0 0 $X=357990 $Y=280205
X377 3 4 ICV_40 $T=358280 358840 1 0 $X=357990 $Y=354630
X378 3 4 ICV_40 $T=366120 280440 0 0 $X=365830 $Y=280205
X379 3 4 ICV_40 $T=398600 327480 0 0 $X=398310 $Y=327245
X380 3 4 ICV_40 $T=399720 249080 1 0 $X=399430 $Y=244870
X381 3 4 ICV_40 $T=400280 264760 0 0 $X=399990 $Y=264525
X382 3 4 ICV_40 $T=408120 264760 0 0 $X=407830 $Y=264525
X383 3 4 ICV_40 $T=408120 303960 0 0 $X=407830 $Y=303725
X384 3 4 ICV_40 $T=417080 241240 0 0 $X=416790 $Y=241005
X385 3 4 ICV_40 $T=419320 303960 0 0 $X=419030 $Y=303725
X386 3 4 ICV_40 $T=433880 272600 0 0 $X=433590 $Y=272365
X387 3 4 ICV_40 $T=440600 303960 0 0 $X=440310 $Y=303725
X388 3 4 ICV_40 $T=442280 335320 1 0 $X=441990 $Y=331110
X389 249 4 255 6 3 NR2D1BWP7T $T=156120 303960 0 0 $X=155830 $Y=303725
X390 253 4 254 250 3 NR2D1BWP7T $T=158360 335320 1 180 $X=155830 $Y=335085
X391 268 4 8 11 3 NR2D1BWP7T $T=160600 351000 0 180 $X=158070 $Y=346790
X392 264 4 266 6 3 NR2D1BWP7T $T=158920 319640 1 0 $X=158630 $Y=315430
X393 249 4 271 265 3 NR2D1BWP7T $T=159480 288280 0 0 $X=159190 $Y=288045
X394 253 4 267 6 3 NR2D1BWP7T $T=161720 327480 1 180 $X=159190 $Y=327245
X395 253 4 269 265 3 NR2D1BWP7T $T=161720 335320 0 180 $X=159190 $Y=331110
X396 13 4 261 11 3 NR2D1BWP7T $T=162280 280440 0 180 $X=159750 $Y=276230
X397 273 4 14 11 3 NR2D1BWP7T $T=162840 358840 0 180 $X=160310 $Y=354630
X398 264 4 274 250 3 NR2D1BWP7T $T=161720 327480 0 0 $X=161430 $Y=327245
X399 264 4 276 265 3 NR2D1BWP7T $T=162280 319640 1 0 $X=161990 $Y=315430
X400 249 4 279 250 3 NR2D1BWP7T $T=164520 343160 1 0 $X=164230 $Y=338950
X401 265 4 283 18 3 NR2D1BWP7T $T=167320 335320 0 0 $X=167030 $Y=335085
X402 284 4 295 18 3 NR2D1BWP7T $T=169000 343160 1 0 $X=168710 $Y=338950
X403 284 4 294 273 3 NR2D1BWP7T $T=169000 343160 0 0 $X=168710 $Y=342925
X404 265 4 286 268 3 NR2D1BWP7T $T=169560 327480 1 0 $X=169270 $Y=323270
X405 253 4 21 11 3 NR2D1BWP7T $T=171800 335320 0 180 $X=169270 $Y=331110
X406 264 4 22 11 3 NR2D1BWP7T $T=172360 327480 1 180 $X=169830 $Y=327245
X407 23 4 285 11 3 NR2D1BWP7T $T=172920 241240 1 180 $X=170390 $Y=241005
X408 273 4 24 258 3 NR2D1BWP7T $T=171800 351000 0 0 $X=171510 $Y=350765
X409 264 4 277 258 3 NR2D1BWP7T $T=175720 288280 0 180 $X=173190 $Y=284070
X410 284 4 296 268 3 NR2D1BWP7T $T=176840 327480 1 180 $X=174310 $Y=327245
X411 30 4 297 31 3 NR2D1BWP7T $T=175160 241240 0 0 $X=174870 $Y=241005
X412 30 4 301 11 3 NR2D1BWP7T $T=179640 241240 1 180 $X=177110 $Y=241005
X413 284 4 289 253 3 NR2D1BWP7T $T=180200 288280 1 180 $X=177670 $Y=288045
X414 284 4 306 264 3 NR2D1BWP7T $T=181320 280440 1 180 $X=178790 $Y=280205
X415 268 4 307 6 3 NR2D1BWP7T $T=184680 335320 1 0 $X=184390 $Y=331110
X416 39 4 323 325 3 NR2D1BWP7T $T=189160 241240 0 0 $X=188870 $Y=241005
X417 325 4 353 56 3 NR2D1BWP7T $T=223880 272600 0 180 $X=221350 $Y=268390
X418 70 4 369 68 3 NR2D1BWP7T $T=234520 327480 0 180 $X=231990 $Y=323270
X419 249 4 352 284 3 NR2D1BWP7T $T=246840 280440 1 180 $X=244310 $Y=280205
X420 88 4 387 11 3 NR2D1BWP7T $T=259720 351000 0 180 $X=257190 $Y=346790
X421 93 4 381 11 3 NR2D1BWP7T $T=260280 319640 0 180 $X=257750 $Y=315430
X422 94 4 391 11 3 NR2D1BWP7T $T=261960 351000 0 180 $X=259430 $Y=346790
X423 96 4 399 11 3 NR2D1BWP7T $T=268120 351000 0 180 $X=265590 $Y=346790
X424 110 4 383 11 3 NR2D1BWP7T $T=288280 343160 1 180 $X=285750 $Y=342925
X425 114 4 113 11 3 NR2D1BWP7T $T=295000 272600 1 180 $X=292470 $Y=272365
X426 70 4 431 115 3 NR2D1BWP7T $T=293320 303960 0 0 $X=293030 $Y=303725
X427 122 4 426 11 3 NR2D1BWP7T $T=296680 280440 0 180 $X=294150 $Y=276230
X428 68 4 435 11 3 NR2D1BWP7T $T=297240 264760 0 180 $X=294710 $Y=260550
X429 121 4 442 123 3 NR2D1BWP7T $T=300040 288280 1 0 $X=299750 $Y=284070
X430 121 4 439 70 3 NR2D1BWP7T $T=304520 335320 1 0 $X=304230 $Y=331110
X431 139 4 444 457 3 NR2D1BWP7T $T=317960 319640 0 180 $X=315430 $Y=315430
X432 102 4 462 115 3 NR2D1BWP7T $T=318520 335320 0 180 $X=315990 $Y=331110
X433 141 4 411 11 3 NR2D1BWP7T $T=326920 241240 1 180 $X=324390 $Y=241005
X434 139 4 464 115 3 NR2D1BWP7T $T=326920 280440 1 180 $X=324390 $Y=280205
X435 123 4 468 457 3 NR2D1BWP7T $T=326920 311800 0 180 $X=324390 $Y=307590
X436 115 4 471 123 3 NR2D1BWP7T $T=324680 343160 0 0 $X=324390 $Y=342925
X437 115 4 425 11 3 NR2D1BWP7T $T=329160 272600 0 180 $X=326630 $Y=268390
X438 121 4 475 148 3 NR2D1BWP7T $T=326920 280440 0 0 $X=326630 $Y=280205
X439 70 4 474 476 3 NR2D1BWP7T $T=328600 335320 1 0 $X=328310 $Y=331110
X440 123 4 477 68 3 NR2D1BWP7T $T=329720 327480 0 0 $X=329430 $Y=327245
X441 121 4 441 139 3 NR2D1BWP7T $T=338680 351000 1 0 $X=338390 $Y=346790
X442 159 4 158 133 3 NR2D1BWP7T $T=346520 256920 1 180 $X=343990 $Y=256685
X443 139 4 456 68 3 NR2D1BWP7T $T=346520 272600 0 180 $X=343990 $Y=268390
X444 70 4 423 457 3 NR2D1BWP7T $T=344280 303960 0 0 $X=343990 $Y=303725
X445 102 4 452 68 3 NR2D1BWP7T $T=347080 264760 1 180 $X=344550 $Y=264525
X446 148 4 488 457 3 NR2D1BWP7T $T=353800 303960 1 180 $X=351270 $Y=303725
X447 102 4 490 476 3 NR2D1BWP7T $T=355480 264760 0 0 $X=355190 $Y=264525
X448 476 4 497 11 3 NR2D1BWP7T $T=358280 256920 1 180 $X=355750 $Y=256685
X449 139 4 495 476 3 NR2D1BWP7T $T=357160 272600 1 0 $X=356870 $Y=268390
X450 121 4 489 172 3 NR2D1BWP7T $T=357160 296120 0 0 $X=356870 $Y=295885
X451 102 4 503 173 3 NR2D1BWP7T $T=357720 264760 0 0 $X=357430 $Y=264525
X452 173 4 498 139 3 NR2D1BWP7T $T=358280 280440 1 0 $X=357990 $Y=276230
X453 172 4 510 457 3 NR2D1BWP7T $T=360520 311800 0 180 $X=357990 $Y=307590
X454 4 3 DCAP64BWP7T $T=408120 296120 0 0 $X=407830 $Y=295885
X492 3 4 ICV_47 $T=156120 264760 1 0 $X=155830 $Y=260550
X493 3 4 ICV_47 $T=198120 249080 1 0 $X=197830 $Y=244870
X494 3 4 ICV_47 $T=198120 288280 0 0 $X=197830 $Y=288045
X495 3 4 ICV_47 $T=198120 311800 0 0 $X=197830 $Y=311565
X496 3 4 ICV_47 $T=198120 319640 1 0 $X=197830 $Y=315430
X497 3 4 ICV_47 $T=198120 358840 1 0 $X=197830 $Y=354630
X498 3 4 ICV_47 $T=240120 264760 1 0 $X=239830 $Y=260550
X499 3 4 ICV_47 $T=282120 249080 1 0 $X=281830 $Y=244870
X500 3 4 ICV_47 $T=282120 311800 0 0 $X=281830 $Y=311565
X501 3 4 ICV_47 $T=282120 327480 0 0 $X=281830 $Y=327245
X502 3 4 ICV_47 $T=282120 358840 1 0 $X=281830 $Y=354630
X503 3 4 ICV_47 $T=324120 249080 0 0 $X=323830 $Y=248845
X504 3 4 ICV_47 $T=324120 264760 1 0 $X=323830 $Y=260550
X505 3 4 ICV_47 $T=324120 272600 0 0 $X=323830 $Y=272365
X506 3 4 ICV_47 $T=324120 288280 1 0 $X=323830 $Y=284070
X507 3 4 ICV_47 $T=324120 327480 1 0 $X=323830 $Y=323270
X508 3 4 ICV_47 $T=324120 351000 0 0 $X=323830 $Y=350765
X509 3 4 ICV_47 $T=366120 256920 1 0 $X=365830 $Y=252710
X510 3 4 ICV_47 $T=366120 280440 1 0 $X=365830 $Y=276230
X511 3 4 ICV_47 $T=366120 311800 0 0 $X=365830 $Y=311565
X512 3 4 ICV_47 $T=366120 335320 0 0 $X=365830 $Y=335085
X513 3 4 ICV_47 $T=366120 343160 1 0 $X=365830 $Y=338950
X514 4 3 DCAP32BWP7T $T=158360 303960 0 0 $X=158070 $Y=303725
X515 4 3 DCAP32BWP7T $T=176840 272600 1 0 $X=176550 $Y=268390
X516 4 3 DCAP32BWP7T $T=178520 351000 0 0 $X=178230 $Y=350765
X517 4 3 DCAP32BWP7T $T=198120 264760 1 0 $X=197830 $Y=260550
X518 4 3 DCAP32BWP7T $T=198120 335320 0 0 $X=197830 $Y=335085
X519 4 3 DCAP32BWP7T $T=198120 351000 1 0 $X=197830 $Y=346790
X520 4 3 DCAP32BWP7T $T=213800 280440 1 0 $X=213510 $Y=276230
X521 4 3 DCAP32BWP7T $T=218840 296120 1 0 $X=218550 $Y=291910
X522 4 3 DCAP32BWP7T $T=221080 335320 1 0 $X=220790 $Y=331110
X523 4 3 DCAP32BWP7T $T=221080 343160 1 0 $X=220790 $Y=338950
X524 4 3 DCAP32BWP7T $T=240120 280440 1 0 $X=239830 $Y=276230
X525 4 3 DCAP32BWP7T $T=240120 303960 1 0 $X=239830 $Y=299750
X526 4 3 DCAP32BWP7T $T=240120 327480 0 0 $X=239830 $Y=327245
X527 4 3 DCAP32BWP7T $T=258600 327480 1 0 $X=258310 $Y=323270
X528 4 3 DCAP32BWP7T $T=260280 358840 1 0 $X=259990 $Y=354630
X529 4 3 DCAP32BWP7T $T=282120 296120 1 0 $X=281830 $Y=291910
X530 4 3 DCAP32BWP7T $T=290520 303960 1 0 $X=290230 $Y=299750
X531 4 3 DCAP32BWP7T $T=293320 264760 0 0 $X=293030 $Y=264525
X532 4 3 DCAP32BWP7T $T=297240 264760 1 0 $X=296950 $Y=260550
X533 4 3 DCAP32BWP7T $T=302280 288280 1 0 $X=301990 $Y=284070
X534 4 3 DCAP32BWP7T $T=303400 343160 0 0 $X=303110 $Y=342925
X535 4 3 DCAP32BWP7T $T=324120 249080 1 0 $X=323830 $Y=244870
X536 4 3 DCAP32BWP7T $T=324120 311800 0 0 $X=323830 $Y=311565
X537 4 3 DCAP32BWP7T $T=324120 319640 1 0 $X=323830 $Y=315430
X538 4 3 DCAP32BWP7T $T=333080 343160 1 0 $X=332790 $Y=338950
X539 4 3 DCAP32BWP7T $T=366120 288280 1 0 $X=365830 $Y=284070
X540 4 3 DCAP32BWP7T $T=366120 327480 1 0 $X=365830 $Y=323270
X541 4 3 DCAP32BWP7T $T=384600 351000 1 0 $X=384310 $Y=346790
X542 4 3 DCAP32BWP7T $T=387400 319640 0 0 $X=387110 $Y=319405
X543 4 3 DCAP32BWP7T $T=408120 280440 1 0 $X=407830 $Y=276230
X544 4 3 DCAP32BWP7T $T=412040 249080 0 0 $X=411750 $Y=248845
X545 4 3 DCAP32BWP7T $T=412040 256920 0 0 $X=411750 $Y=256685
X546 4 3 DCAP32BWP7T $T=415960 272600 0 0 $X=415670 $Y=272365
X547 270 277 289 290 4 3 291 FA1D0BWP7T $T=161160 303960 1 0 $X=160870 $Y=299750
X548 276 296 255 312 4 3 314 FA1D0BWP7T $T=171800 311800 0 0 $X=171510 $Y=311565
X549 295 269 279 317 4 3 318 FA1D0BWP7T $T=175160 343160 1 0 $X=174870 $Y=338950
X550 287 312 302 300 4 3 326 FA1D0BWP7T $T=179640 319640 1 0 $X=179350 $Y=315430
X551 307 283 254 322 4 3 327 FA1D0BWP7T $T=179640 358840 1 0 $X=179350 $Y=354630
X552 351 332 45 44 4 3 42 FA1D0BWP7T $T=211560 241240 1 180 $X=198390 $Y=241005
X553 275 329 298 334 4 3 321 FA1D0BWP7T $T=198680 296120 1 0 $X=198390 $Y=291910
X554 310 267 286 337 4 3 343 FA1D0BWP7T $T=198680 327480 0 0 $X=198390 $Y=327245
X555 294 274 324 338 4 3 49 FA1D0BWP7T $T=198680 343160 0 0 $X=198390 $Y=342925
X556 326 330 339 342 4 3 344 FA1D0BWP7T $T=199800 311800 1 0 $X=199510 $Y=307590
X557 252 304 266 345 4 3 347 FA1D0BWP7T $T=203720 319640 0 0 $X=203430 $Y=319405
X558 320 338 318 335 4 3 333 FA1D0BWP7T $T=221080 335320 0 180 $X=207910 $Y=331110
X559 322 343 54 355 4 3 62 FA1D0BWP7T $T=211000 351000 0 0 $X=210710 $Y=350765
X560 323 297 58 332 4 3 360 FA1D0BWP7T $T=212680 249080 0 0 $X=212390 $Y=248845
X561 317 314 345 339 4 3 368 FA1D0BWP7T $T=218840 319640 0 0 $X=218550 $Y=319405
X562 57 355 333 370 4 3 374 FA1D0BWP7T $T=221640 335320 0 0 $X=221350 $Y=335085
X563 360 359 371 79 4 3 386 FA1D0BWP7T $T=240680 256920 0 0 $X=240390 $Y=256685
X564 335 337 347 380 4 3 379 FA1D0BWP7T $T=240680 319640 0 0 $X=240390 $Y=319405
X565 384 370 379 378 4 3 377 FA1D0BWP7T $T=253560 335320 1 180 $X=240390 $Y=335085
X566 417 401 429 430 4 3 433 FA1D0BWP7T $T=282680 288280 0 0 $X=282390 $Y=288045
X567 432 427 419 416 4 3 417 FA1D0BWP7T $T=295560 319640 1 180 $X=282390 $Y=319405
X568 440 436 421 111 4 3 405 FA1D0BWP7T $T=300600 335320 1 180 $X=287430 $Y=335085
X569 451 444 439 437 4 3 420 FA1D0BWP7T $T=308440 319640 1 180 $X=295270 $Y=319405
X570 422 447 456 449 4 3 458 FA1D0BWP7T $T=302280 311800 1 0 $X=301990 $Y=307590
X571 465 446 449 429 4 3 445 FA1D0BWP7T $T=317400 280440 1 180 $X=304230 $Y=280205
X572 464 442 452 427 4 3 446 FA1D0BWP7T $T=318520 296120 0 180 $X=305350 $Y=291910
X573 484 482 458 470 4 3 467 FA1D0BWP7T $T=337560 296120 0 180 $X=324390 $Y=291910
X574 450 369 471 484 4 3 486 FA1D0BWP7T $T=324680 319640 0 0 $X=324390 $Y=319405
X575 466 483 467 480 4 3 492 FA1D0BWP7T $T=329720 303960 0 0 $X=329430 $Y=303725
X576 475 431 490 465 4 3 494 FA1D0BWP7T $T=331400 280440 0 0 $X=331110 $Y=280205
X577 487 493 499 501 4 3 502 FA1D0BWP7T $T=338120 319640 0 0 $X=337830 $Y=319405
X578 477 157 474 504 4 3 505 FA1D0BWP7T $T=339800 335320 0 0 $X=339510 $Y=335085
X579 489 495 503 496 4 3 493 FA1D0BWP7T $T=340360 296120 1 0 $X=340070 $Y=291910
X580 496 491 494 482 4 3 508 FA1D0BWP7T $T=345400 280440 0 0 $X=345110 $Y=280205
X581 498 164 169 511 4 3 513 FA1D0BWP7T $T=347640 327480 0 0 $X=347350 $Y=327245
X582 519 501 508 483 4 3 518 FA1D0BWP7T $T=379560 303960 1 180 $X=366390 $Y=303725
X583 511 486 504 519 4 3 506 FA1D0BWP7T $T=379560 343160 1 180 $X=366390 $Y=342925
X584 259 3 4 253 INVD1BWP7T $T=158360 327480 0 180 $X=156390 $Y=323270
X585 17 3 4 265 INVD1BWP7T $T=164520 327480 1 0 $X=164230 $Y=323270
X586 280 3 4 249 INVD1BWP7T $T=169000 288280 1 180 $X=167030 $Y=288045
X587 20 3 4 264 INVD1BWP7T $T=169000 280440 1 0 $X=168710 $Y=276230
X588 281 3 4 28 INVD1BWP7T $T=175160 272600 1 0 $X=174870 $Y=268390
X589 305 3 4 32 INVD1BWP7T $T=179640 303960 0 0 $X=179350 $Y=303725
X590 9 3 4 268 INVD1BWP7T $T=186360 327480 1 180 $X=184390 $Y=327245
X591 38 3 4 284 INVD1BWP7T $T=219400 343160 1 0 $X=219110 $Y=338950
X592 356 3 4 31 INVD1BWP7T $T=223320 256920 1 180 $X=221350 $Y=256685
X593 373 3 4 26 INVD1BWP7T $T=257480 343160 0 180 $X=255510 $Y=338950
X594 92 3 4 23 INVD1BWP7T $T=262520 249080 1 180 $X=260550 $Y=248845
X595 103 3 4 418 INVD1BWP7T $T=282680 335320 1 0 $X=282390 $Y=331110
X596 453 3 4 123 INVD1BWP7T $T=315160 327480 1 0 $X=314870 $Y=323270
X597 514 3 4 173 INVD1BWP7T $T=360520 296120 0 180 $X=358550 $Y=291910
X598 500 3 4 148 INVD1BWP7T $T=360520 303960 0 180 $X=358550 $Y=299750
X599 177 3 4 141 INVD1BWP7T $T=368360 249080 1 180 $X=366390 $Y=248845
X600 535 3 4 172 INVD1BWP7T $T=384600 319640 1 180 $X=382630 $Y=319405
X601 174 3 4 476 INVD1BWP7T $T=387400 327480 0 180 $X=385430 $Y=323270
X703 251 3 257 7 4 ND2D1BWP7T $T=156120 343160 0 0 $X=155830 $Y=342925
X704 259 3 278 7 4 ND2D1BWP7T $T=164520 288280 0 0 $X=164230 $Y=288045
X705 280 3 282 7 4 ND2D1BWP7T $T=169000 280440 0 180 $X=166470 $Y=276230
X706 9 3 292 7 4 ND2D1BWP7T $T=172360 327480 0 0 $X=172070 $Y=327245
X707 251 3 27 25 4 ND2D1BWP7T $T=175720 358840 0 180 $X=173190 $Y=354630
X708 259 3 348 41 4 ND2D1BWP7T $T=215480 327480 1 0 $X=215190 $Y=323270
X709 367 3 357 65 4 ND2D1BWP7T $T=232280 249080 1 180 $X=229750 $Y=248845
X710 91 3 87 280 4 ND2D1BWP7T $T=260280 358840 0 180 $X=257750 $Y=354630
X711 92 3 89 65 4 ND2D1BWP7T $T=260840 249080 1 180 $X=258310 $Y=248845
X712 358 3 385 65 4 ND2D1BWP7T $T=273720 272600 0 180 $X=271190 $Y=268390
X713 396 3 108 107 4 ND2D1BWP7T $T=285480 280440 0 180 $X=282950 $Y=276230
X714 367 3 424 389 4 ND2D1BWP7T $T=292760 264760 0 180 $X=290230 $Y=260550
X715 397 3 112 59 4 ND2D1BWP7T $T=292760 272600 1 180 $X=290230 $Y=272365
X716 92 3 438 356 4 ND2D1BWP7T $T=298920 256920 1 180 $X=296390 $Y=256685
X717 120 3 443 363 4 ND2D1BWP7T $T=302280 296120 1 0 $X=301990 $Y=291910
X718 134 3 454 130 4 ND2D1BWP7T $T=311800 335320 1 180 $X=309270 $Y=335085
X719 142 3 472 146 4 ND2D1BWP7T $T=326360 280440 1 0 $X=326070 $Y=276230
X720 146 3 168 138 4 ND2D1BWP7T $T=353800 256920 0 0 $X=353510 $Y=256685
X721 453 3 515 174 4 ND2D1BWP7T $T=358280 303960 0 0 $X=357990 $Y=303725
X722 509 3 516 184 4 ND2D1BWP7T $T=372840 288280 0 0 $X=372550 $Y=288045
X723 514 3 531 448 4 ND2D1BWP7T $T=379000 296120 1 0 $X=378710 $Y=291910
X724 130 3 521 176 4 ND2D1BWP7T $T=394120 351000 0 0 $X=393830 $Y=350765
X725 185 3 530 134 4 ND2D1BWP7T $T=398600 311800 0 180 $X=396070 $Y=307590
X726 160 3 527 532 4 ND2D1BWP7T $T=396360 327480 0 0 $X=396070 $Y=327245
X750 12 3 4 250 INVD0BWP7T $T=160600 351000 0 0 $X=160310 $Y=350765
X751 272 3 4 287 INVD0BWP7T $T=165080 311800 0 0 $X=164790 $Y=311565
X752 290 3 4 298 INVD0BWP7T $T=177960 288280 1 180 $X=175990 $Y=288045
X753 33 3 4 262 INVD0BWP7T $T=181880 303960 0 180 $X=179910 $Y=299750
X754 316 3 4 313 INVD0BWP7T $T=186360 249080 1 180 $X=184390 $Y=248845
X755 299 3 4 330 INVD0BWP7T $T=212120 280440 1 0 $X=211830 $Y=276230
X756 363 3 4 325 INVD0BWP7T $T=233960 272600 1 180 $X=231990 $Y=272365
X757 321 3 4 308 INVD0BWP7T $T=242360 272600 1 180 $X=240390 $Y=272365
X758 416 3 4 413 INVD0BWP7T $T=276520 327480 1 180 $X=274550 $Y=327245
X759 437 3 4 421 INVD0BWP7T $T=286040 335320 0 180 $X=284070 $Y=331110
X760 420 3 4 410 INVD0BWP7T $T=287160 303960 0 180 $X=285190 $Y=299750
X761 460 3 4 432 INVD0BWP7T $T=297240 303960 1 180 $X=295270 $Y=303725
X762 469 3 4 466 INVD0BWP7T $T=326360 280440 0 180 $X=324390 $Y=276230
X763 271 275 16 272 3 4 OAI21D0BWP7T $T=164520 288280 1 180 $X=161430 $Y=288045
X764 352 349 40 316 3 4 OAI21D0BWP7T $T=220520 311800 0 180 $X=217430 $Y=307590
X765 407 402 405 105 3 4 OAI21D0BWP7T $T=271480 311800 0 0 $X=271190 $Y=311565
X766 368 395 380 344 3 4 OAI21D0BWP7T $T=275400 288280 0 180 $X=272310 $Y=284070
X767 408 403 406 105 3 4 OAI21D0BWP7T $T=285480 335320 1 180 $X=282390 $Y=335085
X768 462 440 128 460 3 4 OAI21D0BWP7T $T=318520 311800 0 180 $X=315430 $Y=307590
X769 461 459 433 105 3 4 OAI21D0BWP7T $T=331960 272600 0 180 $X=328870 $Y=268390
X770 172 517 115 516 3 4 OAI21D0BWP7T $T=357720 288280 0 0 $X=357430 $Y=288045
X771 178 522 180 524 3 4 OAI21D0BWP7T $T=370600 264760 0 0 $X=370310 $Y=264525
X772 148 533 68 515 3 4 OAI21D0BWP7T $T=381240 296120 1 0 $X=380950 $Y=291910
X773 178 545 190 536 3 4 OAI21D0BWP7T $T=381800 280440 0 0 $X=381510 $Y=280205
X774 178 525 194 537 3 4 OAI21D0BWP7T $T=388520 264760 0 0 $X=388230 $Y=264525
X775 194 547 195 546 3 4 OAI21D0BWP7T $T=398040 264760 0 180 $X=394950 $Y=260550
X776 178 550 199 549 3 4 OAI21D0BWP7T $T=398600 303960 1 0 $X=398310 $Y=299750
X777 178 541 200 555 3 4 OAI21D0BWP7T $T=398600 311800 1 0 $X=398310 $Y=307590
X778 178 539 201 553 3 4 OAI21D0BWP7T $T=399720 335320 1 0 $X=399430 $Y=331110
X779 190 542 195 554 3 4 OAI21D0BWP7T $T=412040 256920 1 180 $X=408950 $Y=256685
X780 178 543 203 540 3 4 OAI21D0BWP7T $T=413160 319640 0 180 $X=410070 $Y=315430
X781 203 562 195 565 3 4 OAI21D0BWP7T $T=413160 303960 1 0 $X=412870 $Y=299750
X782 204 205 206 207 3 4 OAI21D0BWP7T $T=413720 351000 0 0 $X=413430 $Y=350765
X783 200 558 195 569 3 4 OAI21D0BWP7T $T=416520 303960 0 0 $X=416230 $Y=303725
X784 208 567 210 586 3 4 OAI21D0BWP7T $T=417080 249080 1 0 $X=416790 $Y=244870
X785 201 563 195 568 3 4 OAI21D0BWP7T $T=417640 335320 1 0 $X=417350 $Y=331110
X786 212 560 213 576 3 4 OAI21D0BWP7T $T=422680 343160 1 0 $X=422390 $Y=338950
X787 212 559 206 572 3 4 OAI21D0BWP7T $T=423240 351000 1 0 $X=422950 $Y=346790
X788 208 585 203 574 3 4 OAI21D0BWP7T $T=423800 303960 1 0 $X=423510 $Y=299750
X789 208 566 190 214 3 4 OAI21D0BWP7T $T=427160 256920 0 180 $X=424070 $Y=252710
X790 199 564 195 577 3 4 OAI21D0BWP7T $T=426600 280440 1 0 $X=426310 $Y=276230
X791 208 575 200 578 3 4 OAI21D0BWP7T $T=426600 303960 0 0 $X=426310 $Y=303725
X792 208 584 201 579 3 4 OAI21D0BWP7T $T=433320 335320 0 180 $X=430230 $Y=331110
X793 208 583 194 587 3 4 OAI21D0BWP7T $T=435560 256920 1 180 $X=432470 $Y=256685
X794 213 588 222 591 3 4 OAI21D0BWP7T $T=435000 335320 0 0 $X=434710 $Y=335085
X795 208 580 199 592 3 4 OAI21D0BWP7T $T=436680 264760 1 0 $X=436390 $Y=260550
X796 224 593 222 230 3 4 OAI21D0BWP7T $T=438360 351000 1 0 $X=438070 $Y=346790
X797 231 233 199 238 3 4 OAI21D0BWP7T $T=441160 272600 0 0 $X=440870 $Y=272365
X798 231 589 190 242 3 4 OAI21D0BWP7T $T=441720 256920 1 0 $X=441430 $Y=252710
X799 231 235 203 594 3 4 OAI21D0BWP7T $T=441720 280440 1 0 $X=441430 $Y=276230
X829 16 3 280 17 4 272 ND3D0BWP7T $T=169000 319640 0 180 $X=165910 $Y=315430
X830 40 3 280 38 4 316 ND3D0BWP7T $T=189160 327480 1 180 $X=186070 $Y=327245
X831 63 3 363 65 4 364 ND3D0BWP7T $T=230040 264760 0 0 $X=229750 $Y=264525
X832 128 3 134 136 4 460 ND3D0BWP7T $T=315160 351000 1 0 $X=314870 $Y=346790
X833 170 3 535 130 4 512 ND3D0BWP7T $T=384600 319640 0 0 $X=384310 $Y=319405
X834 3 4 DCAP16BWP7T $T=156120 256920 1 0 $X=155830 $Y=252710
X835 3 4 DCAP16BWP7T $T=158360 343160 0 0 $X=158070 $Y=342925
X836 3 4 DCAP16BWP7T $T=160600 296120 0 0 $X=160310 $Y=295885
X837 3 4 DCAP16BWP7T $T=162840 358840 1 0 $X=162550 $Y=354630
X838 3 4 DCAP16BWP7T $T=169000 319640 1 0 $X=168710 $Y=315430
X839 3 4 DCAP16BWP7T $T=171800 335320 1 0 $X=171510 $Y=331110
X840 3 4 DCAP16BWP7T $T=174040 249080 0 0 $X=173750 $Y=248845
X841 3 4 DCAP16BWP7T $T=179640 241240 0 0 $X=179350 $Y=241005
X842 3 4 DCAP16BWP7T $T=180200 288280 0 0 $X=179910 $Y=288045
X843 3 4 DCAP16BWP7T $T=181320 280440 0 0 $X=181030 $Y=280205
X844 3 4 DCAP16BWP7T $T=181320 296120 0 0 $X=181030 $Y=295885
X845 3 4 DCAP16BWP7T $T=181320 303960 0 0 $X=181030 $Y=303725
X846 3 4 DCAP16BWP7T $T=184680 256920 0 0 $X=184390 $Y=256685
X847 3 4 DCAP16BWP7T $T=184680 311800 0 0 $X=184390 $Y=311565
X848 3 4 DCAP16BWP7T $T=185240 351000 1 0 $X=184950 $Y=346790
X849 3 4 DCAP16BWP7T $T=186360 249080 0 0 $X=186070 $Y=248845
X850 3 4 DCAP16BWP7T $T=186920 272600 0 0 $X=186630 $Y=272365
X851 3 4 DCAP16BWP7T $T=186920 335320 1 0 $X=186630 $Y=331110
X852 3 4 DCAP16BWP7T $T=187480 335320 0 0 $X=187190 $Y=335085
X853 3 4 DCAP16BWP7T $T=198120 296120 0 0 $X=197830 $Y=295885
X854 3 4 DCAP16BWP7T $T=198120 327480 1 0 $X=197830 $Y=323270
X855 3 4 DCAP16BWP7T $T=198120 335320 1 0 $X=197830 $Y=331110
X856 3 4 DCAP16BWP7T $T=198120 351000 0 0 $X=197830 $Y=350765
X857 3 4 DCAP16BWP7T $T=212120 272600 0 0 $X=211830 $Y=272365
X858 3 4 DCAP16BWP7T $T=213240 264760 0 0 $X=212950 $Y=264525
X859 3 4 DCAP16BWP7T $T=216040 256920 1 0 $X=215750 $Y=252710
X860 3 4 DCAP16BWP7T $T=221080 303960 0 0 $X=220790 $Y=303725
X861 3 4 DCAP16BWP7T $T=222760 280440 0 0 $X=222470 $Y=280205
X862 3 4 DCAP16BWP7T $T=229480 241240 0 0 $X=229190 $Y=241005
X863 3 4 DCAP16BWP7T $T=240120 296120 0 0 $X=239830 $Y=295885
X864 3 4 DCAP16BWP7T $T=240120 311800 1 0 $X=239830 $Y=307590
X865 3 4 DCAP16BWP7T $T=240120 327480 1 0 $X=239830 $Y=323270
X866 3 4 DCAP16BWP7T $T=240120 335320 1 0 $X=239830 $Y=331110
X867 3 4 DCAP16BWP7T $T=242360 272600 0 0 $X=242070 $Y=272365
X868 3 4 DCAP16BWP7T $T=253560 335320 0 0 $X=253270 $Y=335085
X869 3 4 DCAP16BWP7T $T=257480 343160 1 0 $X=257190 $Y=338950
X870 3 4 DCAP16BWP7T $T=263080 296120 0 0 $X=262790 $Y=295885
X871 3 4 DCAP16BWP7T $T=263640 288280 1 0 $X=263350 $Y=284070
X872 3 4 DCAP16BWP7T $T=264200 272600 0 0 $X=263910 $Y=272365
X873 3 4 DCAP16BWP7T $T=265320 311800 1 0 $X=265030 $Y=307590
X874 3 4 DCAP16BWP7T $T=271480 343160 1 0 $X=271190 $Y=338950
X875 3 4 DCAP16BWP7T $T=282120 241240 0 0 $X=281830 $Y=241005
X876 3 4 DCAP16BWP7T $T=282120 272600 1 0 $X=281830 $Y=268390
X877 3 4 DCAP16BWP7T $T=282120 280440 0 0 $X=281830 $Y=280205
X878 3 4 DCAP16BWP7T $T=282120 296120 0 0 $X=281830 $Y=295885
X879 3 4 DCAP16BWP7T $T=282120 303960 0 0 $X=281830 $Y=303725
X880 3 4 DCAP16BWP7T $T=282120 351000 0 0 $X=281830 $Y=350765
X881 3 4 DCAP16BWP7T $T=284920 256920 1 0 $X=284630 $Y=252710
X882 3 4 DCAP16BWP7T $T=285480 280440 1 0 $X=285190 $Y=276230
X883 3 4 DCAP16BWP7T $T=311800 335320 0 0 $X=311510 $Y=335085
X884 3 4 DCAP16BWP7T $T=324120 264760 0 0 $X=323830 $Y=264525
X885 3 4 DCAP16BWP7T $T=324120 288280 0 0 $X=323830 $Y=288045
X886 3 4 DCAP16BWP7T $T=334760 256920 0 0 $X=334470 $Y=256685
X887 3 4 DCAP16BWP7T $T=334760 272600 1 0 $X=334470 $Y=268390
X888 3 4 DCAP16BWP7T $T=335320 358840 1 0 $X=335030 $Y=354630
X889 3 4 DCAP16BWP7T $T=337560 343160 0 0 $X=337270 $Y=342925
X890 3 4 DCAP16BWP7T $T=346520 272600 1 0 $X=346230 $Y=268390
X891 3 4 DCAP16BWP7T $T=346520 280440 1 0 $X=346230 $Y=276230
X892 3 4 DCAP16BWP7T $T=349320 256920 1 0 $X=349030 $Y=252710
X893 3 4 DCAP16BWP7T $T=352680 335320 0 0 $X=352390 $Y=335085
X894 3 4 DCAP16BWP7T $T=366120 296120 1 0 $X=365830 $Y=291910
X895 3 4 DCAP16BWP7T $T=366120 319640 0 0 $X=365830 $Y=319405
X896 3 4 DCAP16BWP7T $T=384040 311800 1 0 $X=383750 $Y=307590
X897 3 4 DCAP16BWP7T $T=387400 327480 1 0 $X=387110 $Y=323270
X898 3 4 DCAP16BWP7T $T=391320 264760 0 0 $X=391030 $Y=264525
X899 3 4 DCAP16BWP7T $T=396360 351000 0 0 $X=396070 $Y=350765
X900 3 4 DCAP16BWP7T $T=408120 241240 0 0 $X=407830 $Y=241005
X901 3 4 DCAP16BWP7T $T=408120 288280 0 0 $X=407830 $Y=288045
X902 3 4 DCAP16BWP7T $T=408120 311800 0 0 $X=407830 $Y=311565
X903 3 4 DCAP16BWP7T $T=408120 319640 0 0 $X=407830 $Y=319405
X904 3 4 DCAP16BWP7T $T=408120 335320 1 0 $X=407830 $Y=331110
X905 3 4 DCAP16BWP7T $T=420440 335320 1 0 $X=420150 $Y=331110
X906 3 4 DCAP16BWP7T $T=426040 288280 1 0 $X=425750 $Y=284070
X907 3 4 DCAP16BWP7T $T=429400 280440 1 0 $X=429110 $Y=276230
X908 3 4 DCAP16BWP7T $T=429400 351000 1 0 $X=429110 $Y=346790
X909 3 4 DCAP16BWP7T $T=433320 335320 1 0 $X=433030 $Y=331110
X910 3 4 DCAP16BWP7T $T=437240 311800 1 0 $X=436950 $Y=307590
X911 3 4 DCAP16BWP7T $T=438360 327480 1 0 $X=438070 $Y=323270
X912 3 4 DCAP16BWP7T $T=439480 272600 1 0 $X=439190 $Y=268390
X953 258 3 253 262 252 4 NR3D1BWP7T $T=160600 296120 1 180 $X=155830 $Y=295885
X954 258 3 249 28 270 4 NR3D1BWP7T $T=176280 288280 1 180 $X=171510 $Y=288045
X955 258 3 18 26 29 4 NR3D1BWP7T $T=174040 351000 0 0 $X=173750 $Y=350765
X956 56 3 64 47 359 4 NR3D1BWP7T $T=228920 256920 1 0 $X=228630 $Y=252710
X957 457 3 102 418 451 4 NR3D1BWP7T $T=311800 335320 1 0 $X=311510 $Y=331110
X958 308 300 3 4 291 299 MAOI222D1BWP7T $T=181320 296120 1 180 $X=176550 $Y=295885
X959 313 306 3 4 293 329 MAOI222D1BWP7T $T=198680 272600 0 0 $X=198390 $Y=272365
X960 124 441 3 4 406 436 MAOI222D1BWP7T $T=303400 343160 1 180 $X=298630 $Y=342925
X961 433 445 3 4 470 469 MAOI222D1BWP7T $T=339800 264760 0 0 $X=339510 $Y=264525
X962 28 282 3 270 293 4 AOI21D1BWP7T $T=175160 280440 0 180 $X=171510 $Y=276230
X963 47 357 3 359 351 4 AOI21D1BWP7T $T=221080 264760 1 0 $X=220790 $Y=260550
X964 418 454 3 451 406 4 AOI21D1BWP7T $T=311800 343160 1 0 $X=311510 $Y=338950
X965 433 461 3 459 463 4 AOI21D1BWP7T $T=318520 264760 1 180 $X=314870 $Y=264525
X966 251 18 4 3 INVD2BWP7T $T=169000 343160 0 180 $X=166470 $Y=338950
X967 448 70 4 3 INVD2BWP7T $T=330840 343160 1 0 $X=330550 $Y=338950
X968 160 121 4 3 INVD2BWP7T $T=345400 351000 0 180 $X=342870 $Y=346790
X969 509 139 4 3 INVD2BWP7T $T=358840 296120 0 180 $X=356310 $Y=291910
X1041 5 261 3 4 263 DFQD0BWP7T $T=156120 256920 0 0 $X=155830 $Y=256685
X1042 5 260 3 4 281 DFQD0BWP7T $T=156120 272600 1 0 $X=155830 $Y=268390
X1043 5 285 3 4 256 DFQD0BWP7T $T=168440 256920 1 0 $X=168150 $Y=252710
X1044 5 301 3 4 288 DFQD0BWP7T $T=213240 264760 1 180 $X=202310 $Y=264525
X1045 5 319 3 4 341 DFQD0BWP7T $T=222760 280440 1 180 $X=211830 $Y=280205
X1046 5 346 3 4 305 DFQD0BWP7T $T=223880 296120 1 180 $X=212950 $Y=295885
X1047 5 340 3 4 373 DFQD0BWP7T $T=223880 288280 1 0 $X=223590 $Y=284070
X1048 5 366 3 4 354 DFQD0BWP7T $T=234520 311800 0 180 $X=223590 $Y=307590
X1049 5 76 3 4 376 DFQD0BWP7T $T=251320 288280 0 180 $X=240390 $Y=284070
X1050 5 383 3 4 392 DFQD0BWP7T $T=251320 311800 1 0 $X=251030 $Y=307590
X1051 5 365 3 4 388 DFQD0BWP7T $T=251880 335320 1 0 $X=251590 $Y=331110
X1052 5 387 3 4 361 DFQD0BWP7T $T=263080 296120 1 180 $X=252150 $Y=295885
X1053 5 391 3 4 356 DFQD0BWP7T $T=263640 288280 0 180 $X=252710 $Y=284070
X1054 5 393 3 4 80 DFQD0BWP7T $T=265880 319640 1 180 $X=254950 $Y=319405
X1055 5 85 3 4 382 DFQD0BWP7T $T=255800 256920 0 0 $X=255510 $Y=256685
X1056 5 100 3 4 95 DFQD0BWP7T $T=275400 288280 1 180 $X=264470 $Y=288045
X1057 5 399 3 4 414 DFQD0BWP7T $T=264760 303960 1 0 $X=264470 $Y=299750
X1058 5 398 3 4 103 DFQD0BWP7T $T=264760 335320 0 0 $X=264470 $Y=335085
X1059 5 411 3 4 358 DFQD0BWP7T $T=276520 249080 1 180 $X=265590 $Y=248845
X1060 5 394 3 4 396 DFQD0BWP7T $T=276520 264760 1 180 $X=265590 $Y=264525
X1061 5 412 3 4 397 DFQD0BWP7T $T=276520 280440 0 180 $X=265590 $Y=276230
X1062 5 425 3 4 106 DFQD0BWP7T $T=293320 264760 1 180 $X=282390 $Y=264525
X1063 5 426 3 4 363 DFQD0BWP7T $T=293880 249080 1 180 $X=282950 $Y=248845
X1064 5 119 3 4 367 DFQD0BWP7T $T=303400 241240 1 180 $X=292470 $Y=241005
X1065 5 117 3 4 128 DFQD0BWP7T $T=296120 351000 0 0 $X=295830 $Y=350765
X1066 5 435 3 4 129 DFQD0BWP7T $T=297240 256920 1 0 $X=296950 $Y=252710
X1067 5 455 3 4 126 DFQD0BWP7T $T=315160 241240 1 180 $X=304230 $Y=241005
X1068 150 149 3 4 140 DFQD0BWP7T $T=335320 358840 0 180 $X=324390 $Y=354630
X1069 150 152 3 4 143 DFQD0BWP7T $T=337560 343160 1 180 $X=326630 $Y=342925
X1070 144 497 3 4 154 DFQD0BWP7T $T=349320 256920 0 180 $X=338390 $Y=252710
X1071 144 156 3 4 163 DFQD0BWP7T $T=340360 241240 0 0 $X=340070 $Y=241005
X1072 144 507 3 4 162 DFQD0BWP7T $T=360520 249080 0 180 $X=349590 $Y=244870
X1073 144 526 3 4 175 DFQD0BWP7T $T=377320 241240 1 180 $X=366390 $Y=241005
X1074 144 186 3 4 528 DFQD0BWP7T $T=376760 249080 0 0 $X=376470 $Y=248845
X1075 150 193 3 4 514 DFQD0BWP7T $T=392440 358840 0 180 $X=381510 $Y=354630
X1076 144 547 3 4 538 DFQD0BWP7T $T=399720 249080 0 180 $X=388790 $Y=244870
X1077 144 542 3 4 552 DFQD0BWP7T $T=389640 272600 0 0 $X=389350 $Y=272365
X1078 150 197 3 4 184 DFQD0BWP7T $T=402520 343160 1 180 $X=391590 $Y=342925
X1079 144 558 3 4 557 DFQD0BWP7T $T=408680 311800 1 0 $X=408390 $Y=307590
X1080 150 559 3 4 209 DFQD0BWP7T $T=408680 351000 1 0 $X=408390 $Y=346790
X1081 150 560 3 4 211 DFQD0BWP7T $T=409240 335320 0 0 $X=408950 $Y=335085
X1082 144 562 3 4 544 DFQD0BWP7T $T=409800 296120 1 0 $X=409510 $Y=291910
X1083 150 563 3 4 556 DFQD0BWP7T $T=409800 327480 1 0 $X=409510 $Y=323270
X1084 144 564 3 4 551 DFQD0BWP7T $T=413160 280440 0 0 $X=412870 $Y=280205
X1085 144 567 3 4 561 DFQD0BWP7T $T=424360 256920 0 180 $X=413430 $Y=252710
X1086 144 566 3 4 215 DFQD0BWP7T $T=415400 264760 0 0 $X=415110 $Y=264525
X1087 144 583 3 4 548 DFQD0BWP7T $T=434440 241240 1 180 $X=423510 $Y=241005
X1088 144 585 3 4 570 DFQD0BWP7T $T=435560 296120 0 180 $X=424630 $Y=291910
X1089 150 584 3 4 571 DFQD0BWP7T $T=436120 319640 1 180 $X=425190 $Y=319405
X1090 144 580 3 4 582 DFQD0BWP7T $T=427160 280440 0 0 $X=426870 $Y=280205
X1091 144 589 3 4 216 DFQD0BWP7T $T=439480 272600 0 180 $X=428550 $Y=268390
X1092 150 575 3 4 573 DFQD0BWP7T $T=440600 303960 1 180 $X=429670 $Y=303725
X1093 150 588 3 4 581 DFQD0BWP7T $T=432200 343160 0 0 $X=431910 $Y=342925
X1094 150 593 3 4 218 DFQD0BWP7T $T=442840 358840 0 180 $X=431910 $Y=354630
X1095 32 3 4 268 258 310 NR3D0BWP7T $T=184680 327480 1 180 $X=181590 $Y=327245
X1096 278 302 262 252 3 4 AOI21D0BWP7T $T=177400 303960 1 0 $X=177110 $Y=299750
X1097 292 303 32 310 3 4 AOI21D0BWP7T $T=179640 327480 1 0 $X=179350 $Y=323270
X1098 282 309 28 270 3 4 AOI21D0BWP7T $T=180760 280440 1 0 $X=180470 $Y=276230
X1099 257 320 26 29 3 4 AOI21D0BWP7T $T=189720 343160 1 0 $X=189430 $Y=338950
X1100 407 404 405 402 3 4 AOI21D0BWP7T $T=271480 311800 1 180 $X=268390 $Y=311565
X1101 408 400 406 403 3 4 AOI21D0BWP7T $T=271480 343160 0 180 $X=268390 $Y=338950
X1102 303 3 4 304 BUFFD0BWP7T $T=177400 327480 1 0 $X=177110 $Y=323270
X1103 41 280 3 4 324 AN2D1BWP7T $T=189720 343160 0 0 $X=189430 $Y=342925
X1104 41 20 3 4 52 AN2D1BWP7T $T=216600 343160 1 0 $X=216310 $Y=338950
X1105 358 59 3 4 55 AN2D1BWP7T $T=223880 272600 1 180 $X=220790 $Y=272365
X1106 358 69 3 4 365 AN2D1BWP7T $T=234520 303960 1 180 $X=231430 $Y=303725
X1107 84 280 3 4 82 AN2D1BWP7T $T=258040 358840 0 180 $X=254950 $Y=354630
X1108 97 69 3 4 394 AN2D1BWP7T $T=268680 351000 1 180 $X=265590 $Y=350765
X1109 397 69 3 4 393 AN2D1BWP7T $T=276520 296120 1 180 $X=273430 $Y=295885
X1110 95 107 3 4 109 AN2D1BWP7T $T=288280 272600 1 180 $X=285190 $Y=272365
X1111 430 105 3 4 434 AN2D1BWP7T $T=302840 280440 1 180 $X=299750 $Y=280205
X1112 138 69 3 4 412 AN2D1BWP7T $T=318520 272600 0 180 $X=315430 $Y=268390
X1113 480 105 3 4 481 AN2D1BWP7T $T=331960 272600 1 0 $X=331670 $Y=268390
X1114 184 69 3 4 507 AN2D1BWP7T $T=376200 280440 1 180 $X=373110 $Y=280205
X1115 185 69 3 4 526 AN2D1BWP7T $T=378440 288280 1 180 $X=375350 $Y=288045
X1116 532 69 3 4 188 AN2D1BWP7T $T=384600 351000 0 180 $X=381510 $Y=346790
X1117 300 291 321 4 3 328 XOR3D0BWP7T $T=183000 303960 1 0 $X=182710 $Y=299750
X1118 313 309 306 4 3 315 XNR3D0BWP7T $T=183000 288280 1 0 $X=182710 $Y=284070
X1119 368 344 380 4 3 336 XNR3D0BWP7T $T=251880 303960 1 180 $X=242070 $Y=303725
X1120 37 36 3 315 4 260 35 OAI22D1BWP7T $T=186920 272600 1 180 $X=182710 $Y=272365
X1121 37 43 3 35 4 311 328 OAI22D1BWP7T $T=198680 256920 0 0 $X=198390 $Y=256685
X1122 37 47 3 336 4 340 35 OAI22D1BWP7T $T=212680 256920 1 180 $X=208470 $Y=256685
X1123 368 380 3 384 395 4 IOA21D0BWP7T $T=261960 311800 1 0 $X=261670 $Y=307590
X1124 63 51 378 46 3 4 366 AO22D0BWP7T $T=246840 296120 0 180 $X=242070 $Y=291910
X1125 405 410 413 401 3 4 MAOI222D2BWP7T $T=275960 319640 1 180 $X=268390 $Y=319405
X1126 5 10 3 4 280 DFQD1BWP7T $T=156120 249080 1 0 $X=155830 $Y=244870
X1127 5 34 3 4 251 DFQD1BWP7T $T=180200 256920 1 0 $X=179910 $Y=252710
X1128 5 311 3 4 33 DFQD1BWP7T $T=180200 264760 0 0 $X=179910 $Y=264525
X1129 5 331 3 4 16 DFQD1BWP7T $T=209320 280440 1 180 $X=198390 $Y=280205
X1130 5 350 3 4 40 DFQD1BWP7T $T=234520 296120 1 180 $X=223590 $Y=295885
X1131 5 381 3 4 375 DFQD1BWP7T $T=252440 272600 0 180 $X=241510 $Y=268390
X1132 5 409 3 4 428 DFQD1BWP7T $T=282680 351000 1 0 $X=282390 $Y=346790
X1133 5 404 3 4 415 DFQD1BWP7T $T=289960 311800 1 0 $X=289670 $Y=307590
X1134 5 434 3 4 125 DFQD1BWP7T $T=293320 296120 0 0 $X=293030 $Y=295885
X1135 5 463 3 4 153 DFQD1BWP7T $T=324680 256920 1 0 $X=324390 $Y=252710
X1136 144 473 3 4 485 DFQD1BWP7T $T=326920 241240 0 0 $X=326630 $Y=241005
X1137 5 481 3 4 170 DFQD1BWP7T $T=330840 335320 1 0 $X=330550 $Y=331110
X1138 150 167 3 4 161 DFQD1BWP7T $T=358280 358840 0 180 $X=347350 $Y=354630
X1139 144 182 3 4 509 DFQD1BWP7T $T=377320 256920 1 180 $X=366390 $Y=256685
X1140 144 525 3 4 176 DFQD1BWP7T $T=377320 272600 1 180 $X=366390 $Y=272365
X1141 144 522 3 4 453 DFQD1BWP7T $T=387960 272600 1 180 $X=377030 $Y=272365
X1142 150 539 3 4 532 DFQD1BWP7T $T=391880 343160 1 180 $X=380950 $Y=342925
X1143 150 543 3 4 448 DFQD1BWP7T $T=395240 319640 0 180 $X=384310 $Y=315430
X1144 150 541 3 4 535 DFQD1BWP7T $T=395240 335320 0 180 $X=384310 $Y=331110
X1145 144 550 3 4 500 DFQD1BWP7T $T=402520 296120 1 180 $X=391590 $Y=295885
X1146 46 48 3 4 334 331 35 MOAI22D0BWP7T $T=212120 272600 1 180 $X=207910 $Y=272365
X1147 51 342 3 4 37 346 50 MOAI22D0BWP7T $T=218840 296120 0 180 $X=214630 $Y=291910
X1148 46 53 3 4 35 350 349 MOAI22D0BWP7T $T=221080 303960 1 180 $X=216870 $Y=303725
X1149 46 382 3 4 35 81 362 MOAI22D0BWP7T $T=258600 343160 1 180 $X=254390 $Y=342925
X1150 104 415 3 4 101 99 98 MOAI22D0BWP7T $T=275400 351000 1 180 $X=271190 $Y=350765
X1151 60 348 362 66 372 3 4 XNR4D0BWP7T $T=221640 351000 1 0 $X=221350 $Y=346790
X1152 364 385 90 390 386 3 4 XNR4D0BWP7T $T=251320 272600 0 0 $X=251030 $Y=272365
X1153 529 512 179 521 492 3 4 XNR4D0BWP7T $T=379560 319640 0 180 $X=366390 $Y=315430
X1154 530 527 523 518 505 3 4 XNR4D0BWP7T $T=380680 335320 0 180 $X=367510 $Y=331110
X1155 523 531 529 534 520 3 4 XNR4D0BWP7T $T=393000 303960 1 180 $X=379830 $Y=303725
X1156 72 327 372 374 377 3 4 XOR4D0BWP7T $T=240680 351000 1 0 $X=240390 $Y=346790
X1157 73 75 77 78 382 3 4 XOR4D0BWP7T $T=241240 249080 1 0 $X=240950 $Y=244870
X1158 118 443 390 438 424 3 4 XOR4D0BWP7T $T=298360 272600 1 0 $X=298070 $Y=268390
X1159 137 135 133 132 127 3 4 XOR4D0BWP7T $T=318520 256920 1 180 $X=305350 $Y=256685
X1160 513 506 165 502 161 3 4 XOR4D0BWP7T $T=360520 343160 1 180 $X=347350 $Y=342925
X1161 15 3 4 273 CKND1BWP7T $T=162280 351000 0 0 $X=161990 $Y=350765
X1162 7 3 4 258 CKND1BWP7T $T=164520 319640 1 0 $X=164230 $Y=315430
X1163 389 3 4 86 CKND1BWP7T $T=260280 256920 0 180 $X=258310 $Y=252710
X1164 367 3 4 64 CKND1BWP7T $T=273160 241240 1 180 $X=271190 $Y=241005
X1165 130 3 4 457 CKND1BWP7T $T=346520 303960 0 0 $X=346230 $Y=303725
X1166 124 441 408 124 3 441 4 IAO22D2BWP7T $T=315160 351000 0 180 $X=308710 $Y=346790
X1167 470 445 461 470 3 445 4 IAO22D2BWP7T $T=355480 264760 1 180 $X=349030 $Y=264525
X1168 428 116 3 4 BUFFD1P5BWP7T $T=293320 351000 1 0 $X=293030 $Y=346790
X1169 485 155 3 4 BUFFD1P5BWP7T $T=337560 241240 0 0 $X=337270 $Y=241005
X1170 136 115 4 3 CKND2BWP7T $T=343160 351000 0 180 $X=340630 $Y=346790
X1171 249 4 11 19 3 NR2D0BWP7T $T=165080 351000 1 0 $X=164790 $Y=346790
X1172 102 4 11 409 3 NR2D0BWP7T $T=273160 351000 0 180 $X=270630 $Y=346790
X1173 121 4 11 455 3 NR2D0BWP7T $T=315720 272600 0 180 $X=313190 $Y=268390
X1174 457 4 11 473 3 NR2D0BWP7T $T=338120 264760 1 180 $X=335590 $Y=264525
X1175 187 191 4 178 3 509 189 AOI22D1BWP7T $T=387400 256920 1 180 $X=383190 $Y=256685
X1176 256 3 4 9 CKBD1BWP7T $T=156680 311800 1 0 $X=156390 $Y=307590
X1177 263 3 4 259 CKBD1BWP7T $T=158360 288280 1 0 $X=158070 $Y=284070
X1178 288 3 4 20 CKBD1BWP7T $T=170680 264760 0 0 $X=170390 $Y=264525
X1179 341 3 4 15 CKBD1BWP7T $T=209880 280440 0 0 $X=209590 $Y=280205
X1180 354 3 4 61 CKBD1BWP7T $T=221640 311800 1 0 $X=221350 $Y=307590
X1181 361 3 4 59 CKBD1BWP7T $T=226680 272600 0 0 $X=226390 $Y=272365
X1182 376 3 4 74 CKBD1BWP7T $T=240680 288280 0 0 $X=240390 $Y=288045
X1183 388 3 4 83 CKBD1BWP7T $T=258600 327480 0 180 $X=256070 $Y=323270
X1184 414 3 4 389 CKBD1BWP7T $T=284920 256920 0 180 $X=282390 $Y=252710
X1185 392 3 4 120 CKBD1BWP7T $T=302280 296120 0 180 $X=299750 $Y=291910
X1186 183 3 4 181 CKBD1BWP7T $T=375640 358840 0 180 $X=373110 $Y=354630
X1187 115 516 520 172 517 3 4 OAI31D1BWP7T $T=372840 288280 1 180 $X=368630 $Y=288045
X1188 68 515 534 148 533 3 4 OAI31D1BWP7T $T=388520 327480 1 180 $X=384310 $Y=327245
X1189 63 353 364 4 3 371 OA21D0BWP7T $T=229480 264760 1 0 $X=229190 $Y=260550
X1190 170 510 512 4 3 499 OA21D0BWP7T $T=357160 311800 0 0 $X=356870 $Y=311565
X1191 413 407 416 420 410 4 3 AOI22D0BWP7T $T=282680 311800 1 0 $X=282390 $Y=307590
X1192 528 524 453 187 178 4 3 AOI22D0BWP7T $T=378440 264760 0 0 $X=378150 $Y=264525
X1193 538 537 176 187 178 4 3 AOI22D0BWP7T $T=387960 264760 1 180 $X=384310 $Y=264525
X1194 544 540 448 192 178 4 3 AOI22D0BWP7T $T=389640 296120 0 180 $X=385990 $Y=291910
X1195 195 546 187 538 548 4 3 AOI22D0BWP7T $T=394120 256920 0 0 $X=393830 $Y=256685
X1196 195 196 187 528 198 4 3 AOI22D0BWP7T $T=395800 249080 0 0 $X=395510 $Y=248845
X1197 551 549 500 187 178 4 3 AOI22D0BWP7T $T=399720 272600 0 180 $X=396070 $Y=268390
X1198 556 553 532 192 178 4 3 AOI22D0BWP7T $T=400840 319640 0 180 $X=397190 $Y=315430
X1199 557 555 535 192 178 4 3 AOI22D0BWP7T $T=401400 327480 0 180 $X=397750 $Y=323270
X1200 195 554 187 552 215 4 3 AOI22D0BWP7T $T=399160 264760 1 0 $X=398870 $Y=260550
X1201 552 536 134 187 178 4 3 AOI22D0BWP7T $T=399160 288280 1 0 $X=398870 $Y=284070
X1202 195 202 187 191 561 4 3 AOI22D0BWP7T $T=408680 249080 0 0 $X=408390 $Y=248845
X1203 195 565 192 544 570 4 3 AOI22D0BWP7T $T=417080 288280 0 0 $X=416790 $Y=288045
X1204 195 568 192 556 571 4 3 AOI22D0BWP7T $T=417640 319640 0 0 $X=417350 $Y=319405
X1205 195 569 192 557 573 4 3 AOI22D0BWP7T $T=423240 311800 0 0 $X=422950 $Y=311565
X1206 212 572 192 209 219 4 3 AOI22D0BWP7T $T=426040 351000 1 0 $X=425750 $Y=346790
X1207 212 576 192 211 581 4 3 AOI22D0BWP7T $T=426600 335320 0 0 $X=426310 $Y=335085
X1208 195 577 187 551 582 4 3 AOI22D0BWP7T $T=427160 264760 1 0 $X=426870 $Y=260550
X1209 208 579 192 571 217 4 3 AOI22D0BWP7T $T=427720 327480 0 0 $X=427430 $Y=327245
X1210 208 586 187 561 220 4 3 AOI22D0BWP7T $T=432200 249080 0 0 $X=431910 $Y=248845
X1211 208 574 187 570 239 4 3 AOI22D0BWP7T $T=432200 288280 0 0 $X=431910 $Y=288045
X1212 208 578 187 573 221 4 3 AOI22D0BWP7T $T=432200 311800 0 0 $X=431910 $Y=311565
X1213 208 587 187 548 223 4 3 AOI22D0BWP7T $T=434440 256920 1 0 $X=434150 $Y=252710
X1214 208 592 187 582 240 4 3 AOI22D0BWP7T $T=441160 264760 1 0 $X=440870 $Y=260550
X1215 231 594 237 239 244 4 3 AOI22D0BWP7T $T=441160 296120 1 0 $X=440870 $Y=291910
X1216 222 591 237 581 243 4 3 AOI22D0BWP7T $T=441160 335320 0 0 $X=440870 $Y=335085
X1217 3 4 ICV_76 $T=155000 249080 0 0 $X=154710 $Y=248845
X1218 3 4 ICV_76 $T=155000 280440 0 0 $X=154710 $Y=280205
X1219 3 4 ICV_76 $T=197000 256920 1 0 $X=196710 $Y=252710
X1220 3 4 ICV_76 $T=197000 272600 1 0 $X=196710 $Y=268390
X1221 3 4 ICV_76 $T=197000 288280 1 0 $X=196710 $Y=284070
X1222 3 4 ICV_76 $T=197000 303960 0 0 $X=196710 $Y=303725
X1223 3 4 ICV_76 $T=197000 343160 1 0 $X=196710 $Y=338950
X1224 3 4 ICV_76 $T=239000 249080 0 0 $X=238710 $Y=248845
X1225 3 4 ICV_76 $T=239000 256920 1 0 $X=238710 $Y=252710
X1226 3 4 ICV_76 $T=239000 351000 0 0 $X=238710 $Y=350765
X1227 3 4 ICV_76 $T=281000 288280 1 0 $X=280710 $Y=284070
X1228 3 4 ICV_76 $T=281000 327480 1 0 $X=280710 $Y=323270
X1229 3 4 ICV_76 $T=365000 249080 1 0 $X=364710 $Y=244870
X1230 3 4 ICV_76 $T=365000 272600 1 0 $X=364710 $Y=268390
X1231 3 4 ICV_76 $T=365000 296120 0 0 $X=364710 $Y=295885
X1232 3 4 ICV_76 $T=407000 288280 1 0 $X=406710 $Y=284070
X1233 3 4 ICV_76 $T=407000 327480 0 0 $X=406710 $Y=327245
X1234 3 4 ICV_76 $T=407000 343160 0 0 $X=406710 $Y=342925
X1235 3 4 ICV_76 $T=407000 358840 1 0 $X=406710 $Y=354630
X1236 3 4 ICV_41 $T=156120 241240 0 0 $X=155830 $Y=241005
X1237 3 4 ICV_41 $T=156120 264760 0 0 $X=155830 $Y=264525
X1238 3 4 ICV_41 $T=182440 327480 1 0 $X=182150 $Y=323270
X1239 3 4 ICV_41 $T=183560 280440 1 0 $X=183270 $Y=276230
X1240 3 4 ICV_41 $T=198120 249080 0 0 $X=197830 $Y=248845
X1241 3 4 ICV_41 $T=223320 256920 0 0 $X=223030 $Y=256685
X1242 3 4 ICV_41 $T=223880 351000 0 0 $X=223590 $Y=350765
X1243 3 4 ICV_41 $T=240120 343160 1 0 $X=239830 $Y=338950
X1244 3 4 ICV_41 $T=240120 343160 0 0 $X=239830 $Y=342925
X1245 3 4 ICV_41 $T=240120 358840 1 0 $X=239830 $Y=354630
X1246 3 4 ICV_41 $T=266440 256920 0 0 $X=266150 $Y=256685
X1247 3 4 ICV_41 $T=282120 256920 0 0 $X=281830 $Y=256685
X1248 3 4 ICV_41 $T=307880 256920 1 0 $X=307590 $Y=252710
X1249 3 4 ICV_41 $T=308440 303960 1 0 $X=308150 $Y=299750
X1250 3 4 ICV_41 $T=324120 335320 0 0 $X=323830 $Y=335085
X1251 3 4 ICV_41 $T=324120 351000 1 0 $X=323830 $Y=346790
X1252 3 4 ICV_41 $T=342040 311800 0 0 $X=341750 $Y=311565
X1253 3 4 ICV_41 $T=351000 319640 0 0 $X=350710 $Y=319405
X1254 3 4 ICV_41 $T=351000 343160 1 0 $X=350710 $Y=338950
X1255 3 4 ICV_41 $T=366120 351000 1 0 $X=365830 $Y=346790
X1256 3 4 ICV_41 $T=392440 358840 1 0 $X=392150 $Y=354630
X1257 3 4 ICV_41 $T=393000 303960 0 0 $X=392710 $Y=303725
X1258 3 4 ICV_41 $T=408120 343160 1 0 $X=407830 $Y=338950
X1259 3 4 ICV_41 $T=434440 241240 0 0 $X=434150 $Y=241005
X1260 3 4 ICV_41 $T=434440 351000 0 0 $X=434150 $Y=350765
X1261 3 4 ICV_41 $T=435560 256920 0 0 $X=435270 $Y=256685
X1262 3 4 ICV_37 $T=156120 280440 1 0 $X=155830 $Y=276230
X1263 3 4 ICV_37 $T=156120 288280 0 0 $X=155830 $Y=288045
X1264 3 4 ICV_37 $T=156120 327480 0 0 $X=155830 $Y=327245
X1265 3 4 ICV_37 $T=156120 335320 1 0 $X=155830 $Y=331110
X1266 3 4 ICV_37 $T=165080 256920 1 0 $X=164790 $Y=252710
X1267 3 4 ICV_37 $T=174040 303960 1 0 $X=173750 $Y=299750
X1268 3 4 ICV_37 $T=176280 303960 0 0 $X=175990 $Y=303725
X1269 3 4 ICV_37 $T=184680 249080 1 0 $X=184390 $Y=244870
X1270 3 4 ICV_37 $T=193640 256920 0 0 $X=193350 $Y=256685
X1271 3 4 ICV_37 $T=193640 311800 0 0 $X=193350 $Y=311565
X1272 3 4 ICV_37 $T=207080 351000 0 0 $X=206790 $Y=350765
X1273 3 4 ICV_37 $T=211560 296120 1 0 $X=211270 $Y=291910
X1274 3 4 ICV_37 $T=249080 296120 0 0 $X=248790 $Y=295885
X1275 3 4 ICV_37 $T=262520 264760 0 0 $X=262230 $Y=264525
X1276 3 4 ICV_37 $T=282120 272600 0 0 $X=281830 $Y=272365
X1277 3 4 ICV_37 $T=282120 303960 1 0 $X=281830 $Y=299750
X1278 3 4 ICV_37 $T=293880 256920 1 0 $X=293590 $Y=252710
X1279 3 4 ICV_37 $T=344280 358840 1 0 $X=343990 $Y=354630
X1280 3 4 ICV_37 $T=361640 335320 0 0 $X=361350 $Y=335085
X1281 3 4 ICV_37 $T=380680 335320 1 0 $X=380390 $Y=331110
X1282 3 4 ICV_37 $T=393000 311800 1 0 $X=392710 $Y=307590
X1283 3 4 ICV_37 $T=403640 249080 0 0 $X=403350 $Y=248845
X1284 3 4 ICV_37 $T=436120 319640 0 0 $X=435830 $Y=319405
X1285 3 4 ICV_37 $T=438360 280440 1 0 $X=438070 $Y=276230
X1286 3 4 ICV_60 $T=156120 303960 1 0 $X=155830 $Y=299750
X1287 3 4 ICV_60 $T=174040 280440 0 0 $X=173750 $Y=280205
X1288 3 4 ICV_60 $T=203160 272600 0 0 $X=202870 $Y=272365
X1289 3 4 ICV_60 $T=212680 311800 1 0 $X=212390 $Y=307590
X1290 3 4 ICV_60 $T=224440 264760 1 0 $X=224150 $Y=260550
X1291 3 4 ICV_60 $T=291080 280440 0 0 $X=290790 $Y=280205
X1292 3 4 ICV_60 $T=291080 351000 0 0 $X=290790 $Y=350765
X1293 3 4 ICV_60 $T=333080 288280 0 0 $X=332790 $Y=288045
X1294 3 4 ICV_60 $T=379560 319640 1 0 $X=379270 $Y=315430
X1295 3 4 ICV_60 $T=384040 249080 1 0 $X=383750 $Y=244870
X1296 3 4 ICV_60 $T=408120 280440 0 0 $X=407830 $Y=280205
X1297 3 4 ICV_60 $T=408120 303960 1 0 $X=407830 $Y=299750
X1298 3 4 ICV_60 $T=429960 335320 0 0 $X=429670 $Y=335085
X1299 3 4 ICV_60 $T=443960 264760 0 0 $X=443670 $Y=264525
X1300 3 4 ICV_60 $T=443960 272600 0 0 $X=443670 $Y=272365
X1301 3 4 ICV_60 $T=443960 288280 1 0 $X=443670 $Y=284070
X1302 3 4 ICV_60 $T=443960 296120 0 0 $X=443670 $Y=295885
X1303 3 4 ICV_60 $T=443960 303960 1 0 $X=443670 $Y=299750
X1304 3 4 ICV_43 $T=156120 319640 1 0 $X=155830 $Y=315430
X1305 3 4 ICV_43 $T=169000 288280 0 0 $X=168710 $Y=288045
X1306 3 4 ICV_43 $T=177400 264760 0 0 $X=177110 $Y=264525
X1307 3 4 ICV_43 $T=223880 272600 0 0 $X=223590 $Y=272365
X1308 3 4 ICV_43 $T=249080 335320 1 0 $X=248790 $Y=331110
X1309 3 4 ICV_43 $T=265880 319640 0 0 $X=265590 $Y=319405
X1310 3 4 ICV_43 $T=268680 351000 0 0 $X=268390 $Y=350765
X1311 3 4 ICV_43 $T=309000 343160 1 0 $X=308710 $Y=338950
X1312 3 4 ICV_43 $T=324120 272600 1 0 $X=323830 $Y=268390
X1313 3 4 ICV_43 $T=333080 264760 0 0 $X=332790 $Y=264525
X1314 3 4 ICV_43 $T=337560 296120 1 0 $X=337270 $Y=291910
X1315 3 4 ICV_43 $T=355480 280440 1 0 $X=355190 $Y=276230
X1316 3 4 ICV_43 $T=426040 272600 1 0 $X=425750 $Y=268390
X1317 3 4 ICV_43 $T=429400 288280 0 0 $X=429110 $Y=288045
X1318 3 4 ICV_43 $T=431640 256920 1 0 $X=431350 $Y=252710
X1319 3 4 ICV_43 $T=437800 249080 1 0 $X=437510 $Y=244870
X1320 3 4 ICV_43 $T=446200 311800 1 0 $X=445910 $Y=307590
X1321 3 4 ICV_55 $T=161720 335320 1 0 $X=161430 $Y=331110
X1322 3 4 ICV_55 $T=163960 351000 0 0 $X=163670 $Y=350765
X1323 3 4 ICV_55 $T=189160 288280 0 0 $X=188870 $Y=288045
X1324 3 4 ICV_55 $T=189160 327480 0 0 $X=188870 $Y=327245
X1325 3 4 ICV_55 $T=216040 288280 1 0 $X=215750 $Y=284070
X1326 3 4 ICV_55 $T=222200 264760 0 0 $X=221910 $Y=264525
X1327 3 4 ICV_55 $T=258040 280440 1 0 $X=257750 $Y=276230
X1328 3 4 ICV_55 $T=258040 351000 0 0 $X=257750 $Y=350765
X1329 3 4 ICV_55 $T=273160 241240 0 0 $X=272870 $Y=241005
X1330 3 4 ICV_55 $T=273160 272600 0 0 $X=272870 $Y=272365
X1331 3 4 ICV_55 $T=273160 351000 1 0 $X=272870 $Y=346790
X1332 3 4 ICV_55 $T=315160 264760 1 0 $X=314870 $Y=260550
X1333 3 4 ICV_55 $T=315160 303960 0 0 $X=314870 $Y=303725
X1334 3 4 ICV_55 $T=315160 343160 1 0 $X=314870 $Y=338950
X1335 3 4 ICV_55 $T=342040 249080 1 0 $X=341750 $Y=244870
X1336 3 4 ICV_55 $T=375080 319640 0 0 $X=374790 $Y=319405
X1337 3 4 ICV_55 $T=384040 296120 0 0 $X=383750 $Y=295885
X1338 3 4 ICV_55 $T=388520 327480 0 0 $X=388230 $Y=327245
X1339 3 4 ICV_55 $T=415960 303960 1 0 $X=415670 $Y=299750
X1340 3 4 ICV_55 $T=441160 327480 0 0 $X=440870 $Y=327245
X1341 3 4 ICV_55 $T=441160 351000 1 0 $X=440870 $Y=346790
X1342 3 4 ICV_52 $T=169560 288280 1 0 $X=169270 $Y=284070
X1343 3 4 ICV_52 $T=175720 358840 1 0 $X=175430 $Y=354630
X1344 3 4 ICV_52 $T=180760 335320 1 0 $X=180470 $Y=331110
X1345 3 4 ICV_52 $T=225000 256920 1 0 $X=224710 $Y=252710
X1346 3 4 ICV_52 $T=253560 351000 1 0 $X=253270 $Y=346790
X1347 3 4 ICV_52 $T=260840 288280 0 0 $X=260550 $Y=288045
X1348 3 4 ICV_52 $T=261960 351000 1 0 $X=261670 $Y=346790
X1349 3 4 ICV_52 $T=282120 343160 0 0 $X=281830 $Y=342925
X1350 3 4 ICV_52 $T=286040 311800 1 0 $X=285750 $Y=307590
X1351 3 4 ICV_52 $T=311240 264760 0 0 $X=310950 $Y=264525
X1352 3 4 ICV_52 $T=324120 256920 0 0 $X=323830 $Y=256685
X1353 3 4 ICV_52 $T=372840 249080 0 0 $X=372550 $Y=248845
X1354 3 4 ICV_52 $T=375080 296120 1 0 $X=374790 $Y=291910
X1355 3 4 ICV_52 $T=391880 249080 0 0 $X=391590 $Y=248845
X1356 3 4 ICV_52 $T=403080 296120 1 0 $X=402790 $Y=291910
X1357 3 4 ICV_52 $T=437800 256920 1 0 $X=437510 $Y=252710
X1358 3 4 ICV_54 $T=171800 327480 1 0 $X=171510 $Y=323270
X1359 3 4 ICV_54 $T=175160 280440 1 0 $X=174870 $Y=276230
X1360 3 4 ICV_54 $T=198120 319640 0 0 $X=197830 $Y=319405
X1361 3 4 ICV_54 $T=216040 272600 1 0 $X=215750 $Y=268390
X1362 3 4 ICV_54 $T=216040 335320 0 0 $X=215750 $Y=335085
X1363 3 4 ICV_54 $T=216040 351000 1 0 $X=215750 $Y=346790
X1364 3 4 ICV_54 $T=226680 327480 1 0 $X=226390 $Y=323270
X1365 3 4 ICV_54 $T=233400 256920 1 0 $X=233110 $Y=252710
X1366 3 4 ICV_54 $T=268680 327480 0 0 $X=268390 $Y=327245
X1367 3 4 ICV_54 $T=275400 288280 1 0 $X=275110 $Y=284070
X1368 3 4 ICV_54 $T=275400 288280 0 0 $X=275110 $Y=288045
X1369 3 4 ICV_54 $T=324120 327480 0 0 $X=323830 $Y=327245
X1370 3 4 ICV_54 $T=359400 335320 1 0 $X=359110 $Y=331110
X1371 3 4 ICV_54 $T=376200 280440 0 0 $X=375910 $Y=280205
X1372 3 4 ICV_54 $T=377320 256920 0 0 $X=377030 $Y=256685
X1373 3 4 ICV_54 $T=393000 303960 1 0 $X=392710 $Y=299750
X1374 3 4 ICV_54 $T=401400 303960 1 0 $X=401110 $Y=299750
X1375 3 4 ICV_54 $T=401400 311800 1 0 $X=401110 $Y=307590
X1376 3 4 ICV_54 $T=408120 256920 1 0 $X=407830 $Y=252710
X1377 3 4 ICV_54 $T=408120 351000 0 0 $X=407830 $Y=350765
X1378 3 4 ICV_54 $T=426600 311800 0 0 $X=426310 $Y=311565
X1379 3 4 ICV_54 $T=435560 296120 1 0 $X=435270 $Y=291910
X1380 3 4 ICV_54 $T=443400 311800 0 0 $X=443110 $Y=311565
X1381 3 4 ICV_54 $T=443400 319640 0 0 $X=443110 $Y=319405
X1382 3 4 ICV_54 $T=443400 343160 1 0 $X=443110 $Y=338950
X1383 325 4 11 319 3 NR2XD0BWP7T $T=190840 249080 0 180 $X=188310 $Y=244870
X1384 67 4 11 71 3 NR2XD0BWP7T $T=232280 249080 0 0 $X=231990 $Y=248845
X1385 3 4 ICV_38 $T=192520 319640 1 0 $X=192230 $Y=315430
X1386 3 4 ICV_38 $T=192520 358840 1 0 $X=192230 $Y=354630
X1387 3 4 ICV_38 $T=234520 296120 0 0 $X=234230 $Y=295885
X1388 3 4 ICV_38 $T=234520 303960 0 0 $X=234230 $Y=303725
X1389 3 4 ICV_38 $T=234520 311800 1 0 $X=234230 $Y=307590
X1390 3 4 ICV_38 $T=234520 327480 1 0 $X=234230 $Y=323270
X1391 3 4 ICV_38 $T=276520 249080 0 0 $X=276230 $Y=248845
X1392 3 4 ICV_38 $T=276520 280440 1 0 $X=276230 $Y=276230
X1393 3 4 ICV_38 $T=276520 296120 0 0 $X=276230 $Y=295885
X1394 3 4 ICV_38 $T=276520 327480 0 0 $X=276230 $Y=327245
X1395 3 4 ICV_38 $T=276520 343160 0 0 $X=276230 $Y=342925
X1396 3 4 ICV_38 $T=318520 256920 0 0 $X=318230 $Y=256685
X1397 3 4 ICV_38 $T=318520 264760 0 0 $X=318230 $Y=264525
X1398 3 4 ICV_38 $T=318520 272600 1 0 $X=318230 $Y=268390
X1399 3 4 ICV_38 $T=318520 335320 1 0 $X=318230 $Y=331110
X1400 3 4 ICV_38 $T=360520 280440 1 0 $X=360230 $Y=276230
X1401 3 4 ICV_38 $T=360520 296120 1 0 $X=360230 $Y=291910
X1402 3 4 ICV_38 $T=360520 327480 0 0 $X=360230 $Y=327245
X1403 3 4 ICV_38 $T=402520 280440 0 0 $X=402230 $Y=280205
X1404 3 4 ICV_38 $T=402520 296120 0 0 $X=402230 $Y=295885
X1405 3 4 ICV_38 $T=402520 335320 1 0 $X=402230 $Y=331110
X1406 3 4 ICV_45 $T=211560 327480 0 0 $X=211270 $Y=327245
X1407 3 4 ICV_45 $T=211560 343160 0 0 $X=211270 $Y=342925
X1408 3 4 ICV_45 $T=240120 241240 0 0 $X=239830 $Y=241005
X1409 3 4 ICV_45 $T=240120 311800 0 0 $X=239830 $Y=311565
X1410 3 4 ICV_45 $T=246840 280440 0 0 $X=246550 $Y=280205
X1411 3 4 ICV_45 $T=246840 296120 1 0 $X=246550 $Y=291910
X1412 3 4 ICV_45 $T=254120 249080 1 0 $X=253830 $Y=244870
X1413 3 4 ICV_45 $T=282120 319640 1 0 $X=281830 $Y=315430
X1414 3 4 ICV_45 $T=282120 343160 1 0 $X=281830 $Y=338950
X1415 3 4 ICV_45 $T=293880 249080 0 0 $X=293590 $Y=248845
X1416 3 4 ICV_45 $T=295000 272600 0 0 $X=294710 $Y=272365
X1417 3 4 ICV_45 $T=295560 288280 0 0 $X=295270 $Y=288045
X1418 3 4 ICV_45 $T=326920 311800 1 0 $X=326630 $Y=307590
X1419 3 4 ICV_45 $T=366120 264760 1 0 $X=365830 $Y=260550
X1420 3 4 ICV_45 $T=377320 241240 0 0 $X=377030 $Y=241005
X1421 3 4 ICV_45 $T=378440 288280 0 0 $X=378150 $Y=288045
X1422 35 51 3 4 INVD2P5BWP7T $T=219400 264760 0 180 $X=216310 $Y=260550
X1423 375 3 4 65 BUFFD3BWP7T $T=240680 264760 0 0 $X=240390 $Y=264525
X1424 400 3 4 398 BUFFD1BWP7T $T=268680 327480 1 180 $X=266150 $Y=327245
X1425 415 423 3 4 422 419 IAO21D0BWP7T $T=290520 303960 0 180 $X=286870 $Y=299750
X1426 125 468 3 4 450 447 IAO21D0BWP7T $T=324680 303960 0 0 $X=324390 $Y=303725
X1427 153 488 3 4 487 491 IAO21D0BWP7T $T=338120 288280 0 0 $X=337830 $Y=288045
X1428 130 448 415 4 3 422 AN3D1BWP7T $T=307880 335320 1 180 $X=304230 $Y=335085
X1429 130 453 125 4 3 450 AN3D1BWP7T $T=310120 335320 0 180 $X=306470 $Y=331110
X1430 130 500 153 4 3 487 AN3D1BWP7T $T=348200 303960 0 0 $X=347910 $Y=303725
X1431 131 5 3 4 INVD12BWP7T $T=309000 319640 0 0 $X=308710 $Y=319405
X1432 171 4 166 3 CKND12BWP7T $T=357720 319640 0 180 $X=348470 $Y=315430
X1433 144 545 134 3 4 DFQD2BWP7T $T=397480 288280 0 180 $X=385990 $Y=284070
X1434 192 3 4 187 BUFFD5BWP7T $T=415960 272600 1 180 $X=409510 $Y=272365
X1435 590 225 3 4 BUFFD2BWP7T $T=436680 303960 1 0 $X=436390 $Y=299750
X1436 227 178 228 3 4 ND2D2BWP7T $T=441160 327480 1 180 $X=436950 $Y=327245
X1437 228 3 229 208 4 CKND2D2BWP7T $T=443400 311800 1 180 $X=439190 $Y=311565
X1438 226 3 227 590 4 CKND2D2BWP7T $T=440040 303960 1 0 $X=439750 $Y=299750
X1439 236 195 228 3 4 ND2D1P5BWP7T $T=443400 319640 1 180 $X=439190 $Y=319405
X1440 229 232 226 3 4 ND2D1P5BWP7T $T=443960 288280 0 180 $X=439750 $Y=284070
X1441 236 234 241 3 4 ND2D1P5BWP7T $T=444520 249080 0 180 $X=440310 $Y=244870
.ENDS
***************************************
.SUBCKT __$$VIA34_520_520_21_58
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_80 1 2
** N=2 EP=2 IP=4 FDC=48
*.SEEDPROM
X1 2 1 DCAP64BWP7T $T=1120 0 0 0 $X=830 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_64 1 2
** N=2 EP=2 IP=4 FDC=6
*.SEEDPROM
X0 1 2 DCAP8BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_81 1 2
** N=2 EP=2 IP=4 FDC=54
*.SEEDPROM
X0 1 2 ICV_80 $T=0 0 0 0 $X=-290 $Y=-235
X1 1 2 ICV_64 $T=36960 0 0 0 $X=36670 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_69 1 2
** N=2 EP=2 IP=4 FDC=12
*.SEEDPROM
X1 1 2 DCAP16BWP7T $T=1120 0 0 0 $X=830 $Y=-235
.ENDS
***************************************
.SUBCKT OAI211D1BWP7T C VSS B A1 VDD ZN A2
** N=10 EP=7 IP=0 FDC=8
*.SEEDPROM
M0 9 C VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 8 B 9 VSS N L=1.8e-07 W=1e-06 $X=1120 $Y=345 $D=0
M2 ZN A1 8 VSS N L=1.8e-07 W=1e-06 $X=1840 $Y=345 $D=0
M3 8 A2 ZN VSS N L=1.8e-07 W=1e-06 $X=2560 $Y=345 $D=0
M4 ZN C VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M5 VDD B ZN VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M6 10 A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M7 ZN A2 10 VDD P L=1.8e-07 W=1.37e-06 $X=2560 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ND2D4BWP7T A2 VSS A1 ZN VDD
** N=6 EP=5 IP=0 FDC=16
*.SEEDPROM
M0 VSS A2 6 VSS N L=1.8e-07 W=1e-06 $X=720 $Y=345 $D=0
M1 6 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=1440 $Y=345 $D=0
M2 VSS A2 6 VSS N L=1.8e-07 W=1e-06 $X=2160 $Y=345 $D=0
M3 6 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=2880 $Y=345 $D=0
M4 ZN A1 6 VSS N L=1.8e-07 W=1e-06 $X=3600 $Y=345 $D=0
M5 6 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=4325 $Y=345 $D=0
M6 ZN A1 6 VSS N L=1.8e-07 W=1e-06 $X=5045 $Y=345 $D=0
M7 6 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=5765 $Y=345 $D=0
M8 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=720 $Y=2205 $D=16
M9 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1440 $Y=2205 $D=16
M10 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2160 $Y=2205 $D=16
M11 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2880 $Y=2205 $D=16
M12 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3600 $Y=2205 $D=16
M13 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4325 $Y=2205 $D=16
M14 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=5045 $Y=2205 $D=16
M15 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=5765 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR2XD3BWP7T A2 VDD A1 VSS ZN
** N=6 EP=5 IP=0 FDC=20
*.SEEDPROM
M0 VSS A2 ZN VSS N L=1.8e-07 W=6e-07 $X=820 $Y=345 $D=0
M1 ZN A2 VSS VSS N L=1.8e-07 W=6e-07 $X=1540 $Y=345 $D=0
M2 VSS A2 ZN VSS N L=1.8e-07 W=6e-07 $X=2260 $Y=345 $D=0
M3 ZN A2 VSS VSS N L=1.8e-07 W=6e-07 $X=2980 $Y=345 $D=0
M4 VSS A2 ZN VSS N L=1.8e-07 W=6e-07 $X=3700 $Y=345 $D=0
M5 ZN A1 VSS VSS N L=1.8e-07 W=6e-07 $X=4420 $Y=345 $D=0
M6 VSS A1 ZN VSS N L=1.8e-07 W=6e-07 $X=5140 $Y=345 $D=0
M7 ZN A1 VSS VSS N L=1.8e-07 W=6e-07 $X=5860 $Y=345 $D=0
M8 VSS A1 ZN VSS N L=1.8e-07 W=6e-07 $X=6580 $Y=345 $D=0
M9 ZN A1 VSS VSS N L=1.8e-07 W=6e-07 $X=7300 $Y=345 $D=0
M10 6 A2 VDD VDD P L=1.8e-07 W=1.14e-06 $X=820 $Y=2435 $D=16
M11 VDD A2 6 VDD P L=1.8e-07 W=1.77e-06 $X=1540 $Y=1805 $D=16
M12 6 A2 VDD VDD P L=1.8e-07 W=1.77e-06 $X=2260 $Y=1805 $D=16
M13 VDD A2 6 VDD P L=1.8e-07 W=1.77e-06 $X=2980 $Y=1805 $D=16
M14 6 A2 VDD VDD P L=1.8e-07 W=1.77e-06 $X=3700 $Y=1805 $D=16
M15 ZN A1 6 VDD P L=1.8e-07 W=1.77e-06 $X=4420 $Y=1805 $D=16
M16 6 A1 ZN VDD P L=1.8e-07 W=1.77e-06 $X=5140 $Y=1805 $D=16
M17 ZN A1 6 VDD P L=1.8e-07 W=1.77e-06 $X=5860 $Y=1805 $D=16
M18 6 A1 ZN VDD P L=1.8e-07 W=1.77e-06 $X=6580 $Y=1805 $D=16
M19 ZN A1 6 VDD P L=1.8e-07 W=1.14e-06 $X=7300 $Y=2435 $D=16
.ENDS
***************************************
.SUBCKT MOAI22D1BWP7T B1 B2 VSS A1 ZN A2 VDD
** N=11 EP=7 IP=0 FDC=10
*.SEEDPROM
M0 10 B1 8 VSS N L=1.8e-07 W=1e-06 $X=705 $Y=345 $D=0
M1 VSS B2 10 VSS N L=1.8e-07 W=1e-06 $X=1265 $Y=345 $D=0
M2 9 8 VSS VSS N L=1.8e-07 W=1e-06 $X=2025 $Y=345 $D=0
M3 ZN A1 9 VSS N L=1.8e-07 W=1e-06 $X=2745 $Y=345 $D=0
M4 9 A2 ZN VSS N L=1.8e-07 W=1e-06 $X=3465 $Y=345 $D=0
M5 8 B1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=705 $Y=2205 $D=16
M6 VDD B2 8 VDD P L=1.8e-07 W=1.37e-06 $X=1425 $Y=2205 $D=16
M7 ZN 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2265 $Y=2205 $D=16
M8 11 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2985 $Y=2205 $D=16
M9 VDD A2 11 VDD P L=1.8e-07 W=1.37e-06 $X=3585 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AOI211D1BWP7T C VDD B A2 VSS ZN A1
** N=10 EP=7 IP=0 FDC=8
*.SEEDPROM
M0 ZN C VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS B ZN VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 9 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=2060 $Y=345 $D=0
M3 ZN A1 9 VSS N L=1.8e-07 W=1e-06 $X=2560 $Y=345 $D=0
M4 10 C VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M5 8 B 10 VDD P L=1.8e-07 W=1.37e-06 $X=1120 $Y=2205 $D=16
M6 ZN A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=1840 $Y=2205 $D=16
M7 8 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2560 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR2D1P5BWP7T A1 ZN A2 VDD VSS
** N=7 EP=5 IP=0 FDC=8
*.SEEDPROM
M0 ZN A2 VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS A1 ZN VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 ZN A1 VSS VSS N L=1.8e-07 W=5e-07 $X=2080 $Y=345 $D=0
M3 VSS A2 ZN VSS N L=1.8e-07 W=5e-07 $X=2800 $Y=345 $D=0
M4 6 A2 VDD VDD P L=1.8e-07 W=1.03e-06 $X=620 $Y=2545 $D=16
M5 ZN A1 6 VDD P L=1.8e-07 W=1.03e-06 $X=1220 $Y=2545 $D=16
M6 7 A1 ZN VDD P L=1.8e-07 W=1.03e-06 $X=1940 $Y=2545 $D=16
M7 VDD A2 7 VDD P L=1.8e-07 W=1.03e-06 $X=2800 $Y=2545 $D=16
.ENDS
***************************************
.SUBCKT BUFFD8BWP7T I Z VSS VDD
** N=5 EP=4 IP=0 FDC=22
*.SEEDPROM
M0 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 5 I VSS VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=2060 $Y=345 $D=0
M3 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=2780 $Y=345 $D=0
M4 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=3500 $Y=345 $D=0
M5 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=4220 $Y=345 $D=0
M6 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=4940 $Y=345 $D=0
M7 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=5660 $Y=345 $D=0
M8 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=6380 $Y=345 $D=0
M9 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=7100 $Y=345 $D=0
M10 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=7820 $Y=345 $D=0
M11 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M12 5 I VDD VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M13 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M14 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M15 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=3500 $Y=2205 $D=16
M16 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4220 $Y=2205 $D=16
M17 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=4940 $Y=2205 $D=16
M18 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=5660 $Y=2205 $D=16
M19 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=6380 $Y=2205 $D=16
M20 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=7100 $Y=2205 $D=16
M21 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=7820 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_82 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279
** N=659 EP=278 IP=4620 FDC=11816
*.SEEDPROM
M0 101 97 3 3 N L=1.8e-07 W=1e-06 $X=305800 $Y=476785 $D=0
M1 3 97 101 3 N L=1.8e-07 W=1e-06 $X=306520 $Y=476785 $D=0
M2 101 97 3 3 N L=1.8e-07 W=1e-06 $X=307280 $Y=476785 $D=0
M3 3 97 101 3 N L=1.8e-07 W=1e-06 $X=308000 $Y=476785 $D=0
M4 101 97 3 3 N L=1.8e-07 W=1e-06 $X=308760 $Y=476785 $D=0
M5 101 97 1 1 P L=1.8e-07 W=1.37e-06 $X=305800 $Y=478645 $D=16
M6 1 97 101 1 P L=1.8e-07 W=1.37e-06 $X=306520 $Y=478645 $D=16
M7 101 97 1 1 P L=1.8e-07 W=1.37e-06 $X=307280 $Y=478645 $D=16
M8 1 97 101 1 P L=1.8e-07 W=1.37e-06 $X=308000 $Y=478645 $D=16
M9 101 97 1 1 P L=1.8e-07 W=1.37e-06 $X=308760 $Y=478645 $D=16
X28 4 3 PVSS3CDG $T=0 450000 0 270 $X=0 $Y=369400
X202 1 3 DCAPBWP7T $T=167320 366680 1 0 $X=167030 $Y=362470
X203 1 3 DCAPBWP7T $T=167320 374520 0 0 $X=167030 $Y=374285
X204 1 3 DCAPBWP7T $T=169560 405880 1 0 $X=169270 $Y=401670
X205 1 3 DCAPBWP7T $T=169560 445080 1 0 $X=169270 $Y=440870
X206 1 3 DCAPBWP7T $T=195320 366680 1 0 $X=195030 $Y=362470
X207 1 3 DCAPBWP7T $T=195320 366680 0 0 $X=195030 $Y=366445
X208 1 3 DCAPBWP7T $T=207080 413720 1 0 $X=206790 $Y=409510
X209 1 3 DCAPBWP7T $T=211560 358840 0 0 $X=211270 $Y=358605
X210 1 3 DCAPBWP7T $T=229480 390200 0 0 $X=229190 $Y=389965
X211 1 3 DCAPBWP7T $T=237320 390200 0 0 $X=237030 $Y=389965
X212 1 3 DCAPBWP7T $T=237320 413720 1 0 $X=237030 $Y=409510
X213 1 3 DCAPBWP7T $T=237320 421560 0 0 $X=237030 $Y=421325
X214 1 3 DCAPBWP7T $T=237320 445080 0 0 $X=237030 $Y=444845
X215 1 3 DCAPBWP7T $T=237320 460760 0 0 $X=237030 $Y=460525
X216 1 3 DCAPBWP7T $T=249640 445080 1 0 $X=249350 $Y=440870
X217 1 3 DCAPBWP7T $T=253000 398040 0 0 $X=252710 $Y=397805
X218 1 3 DCAPBWP7T $T=253000 429400 1 0 $X=252710 $Y=425190
X219 1 3 DCAPBWP7T $T=253560 437240 0 0 $X=253270 $Y=437005
X220 1 3 DCAPBWP7T $T=258040 405880 1 0 $X=257750 $Y=401670
X221 1 3 DCAPBWP7T $T=260280 421560 0 0 $X=259990 $Y=421325
X222 1 3 DCAPBWP7T $T=263640 452920 0 0 $X=263350 $Y=452685
X223 1 3 DCAPBWP7T $T=263640 468600 1 0 $X=263350 $Y=464390
X224 1 3 DCAPBWP7T $T=264760 437240 0 0 $X=264470 $Y=437005
X225 1 3 DCAPBWP7T $T=265320 366680 1 0 $X=265030 $Y=362470
X226 1 3 DCAPBWP7T $T=279320 358840 0 0 $X=279030 $Y=358605
X227 1 3 DCAPBWP7T $T=279320 405880 1 0 $X=279030 $Y=401670
X228 1 3 DCAPBWP7T $T=279320 421560 1 0 $X=279030 $Y=417350
X229 1 3 DCAPBWP7T $T=279320 429400 0 0 $X=279030 $Y=429165
X230 1 3 DCAPBWP7T $T=291080 445080 1 0 $X=290790 $Y=440870
X231 1 3 DCAPBWP7T $T=293320 452920 0 0 $X=293030 $Y=452685
X232 1 3 DCAPBWP7T $T=306200 358840 0 0 $X=305910 $Y=358605
X233 1 3 DCAPBWP7T $T=314600 429400 1 0 $X=314310 $Y=425190
X234 1 3 DCAPBWP7T $T=321320 382360 1 0 $X=321030 $Y=378150
X235 1 3 DCAPBWP7T $T=321320 421560 1 0 $X=321030 $Y=417350
X236 1 3 DCAPBWP7T $T=321320 452920 0 0 $X=321030 $Y=452685
X237 1 3 DCAPBWP7T $T=321320 468600 1 0 $X=321030 $Y=464390
X238 1 3 DCAPBWP7T $T=324120 390200 0 0 $X=323830 $Y=389965
X239 1 3 DCAPBWP7T $T=337560 374520 1 0 $X=337270 $Y=370310
X240 1 3 DCAPBWP7T $T=337560 382360 0 0 $X=337270 $Y=382125
X241 1 3 DCAPBWP7T $T=348200 460760 0 0 $X=347910 $Y=460525
X242 1 3 DCAPBWP7T $T=356040 437240 0 0 $X=355750 $Y=437005
X243 1 3 DCAPBWP7T $T=356600 460760 1 0 $X=356310 $Y=456550
X244 1 3 DCAPBWP7T $T=363320 374520 1 0 $X=363030 $Y=370310
X245 1 3 DCAPBWP7T $T=363320 398040 0 0 $X=363030 $Y=397805
X246 1 3 DCAPBWP7T $T=363320 445080 0 0 $X=363030 $Y=444845
X247 1 3 DCAPBWP7T $T=363320 452920 0 0 $X=363030 $Y=452685
X248 1 3 DCAPBWP7T $T=363320 468600 1 0 $X=363030 $Y=464390
X249 1 3 DCAPBWP7T $T=363320 468600 0 0 $X=363030 $Y=468365
X250 1 3 DCAPBWP7T $T=363320 476440 0 0 $X=363030 $Y=476205
X251 1 3 DCAPBWP7T $T=366120 484280 1 0 $X=365830 $Y=480070
X252 1 3 DCAPBWP7T $T=370600 429400 0 0 $X=370310 $Y=429165
X253 1 3 DCAPBWP7T $T=376200 476440 0 0 $X=375910 $Y=476205
X254 1 3 DCAPBWP7T $T=388520 382360 1 0 $X=388230 $Y=378150
X255 1 3 DCAPBWP7T $T=390760 429400 0 0 $X=390470 $Y=429165
X256 1 3 DCAPBWP7T $T=398040 468600 1 0 $X=397750 $Y=464390
X257 1 3 DCAPBWP7T $T=398600 437240 1 0 $X=398310 $Y=433030
X258 1 3 DCAPBWP7T $T=405320 398040 1 0 $X=405030 $Y=393830
X259 1 3 DCAPBWP7T $T=405320 421560 1 0 $X=405030 $Y=417350
X260 1 3 DCAPBWP7T $T=408120 413720 1 0 $X=407830 $Y=409510
X261 1 3 DCAPBWP7T $T=410920 445080 1 0 $X=410630 $Y=440870
X262 1 3 DCAPBWP7T $T=416520 445080 0 0 $X=416230 $Y=444845
X263 1 3 DCAPBWP7T $T=423800 452920 0 0 $X=423510 $Y=452685
X264 1 3 DCAPBWP7T $T=432760 413720 0 0 $X=432470 $Y=413485
X265 1 3 DCAPBWP7T $T=440040 437240 0 0 $X=439750 $Y=437005
X266 1 3 DCAPBWP7T $T=447320 390200 1 0 $X=447030 $Y=385990
X267 1 3 DCAPBWP7T $T=447320 405880 1 0 $X=447030 $Y=401670
X268 1 3 DCAPBWP7T $T=447320 460760 0 0 $X=447030 $Y=460525
X269 3 1 DCAP8BWP7T $T=156120 405880 1 0 $X=155830 $Y=401670
X270 3 1 DCAP8BWP7T $T=156120 445080 1 0 $X=155830 $Y=440870
X271 3 1 DCAP8BWP7T $T=156120 484280 1 0 $X=155830 $Y=480070
X272 3 1 DCAP8BWP7T $T=192520 390200 1 0 $X=192230 $Y=385990
X273 3 1 DCAP8BWP7T $T=192520 421560 1 0 $X=192230 $Y=417350
X274 3 1 DCAP8BWP7T $T=192520 437240 1 0 $X=192230 $Y=433030
X275 3 1 DCAP8BWP7T $T=192520 460760 0 0 $X=192230 $Y=460525
X276 3 1 DCAP8BWP7T $T=198120 390200 1 0 $X=197830 $Y=385990
X277 3 1 DCAP8BWP7T $T=211560 421560 1 0 $X=211270 $Y=417350
X278 3 1 DCAP8BWP7T $T=216040 382360 1 0 $X=215750 $Y=378150
X279 3 1 DCAP8BWP7T $T=216040 398040 1 0 $X=215750 $Y=393830
X280 3 1 DCAP8BWP7T $T=224440 437240 1 0 $X=224150 $Y=433030
X281 3 1 DCAP8BWP7T $T=225000 390200 0 0 $X=224710 $Y=389965
X282 3 1 DCAP8BWP7T $T=232840 390200 0 0 $X=232550 $Y=389965
X283 3 1 DCAP8BWP7T $T=232840 445080 0 0 $X=232550 $Y=444845
X284 3 1 DCAP8BWP7T $T=234520 366680 1 0 $X=234230 $Y=362470
X285 3 1 DCAP8BWP7T $T=234520 405880 0 0 $X=234230 $Y=405645
X286 3 1 DCAP8BWP7T $T=234520 460760 1 0 $X=234230 $Y=456550
X287 3 1 DCAP8BWP7T $T=240120 429400 1 0 $X=239830 $Y=425190
X288 3 1 DCAP8BWP7T $T=240120 484280 1 0 $X=239830 $Y=480070
X289 3 1 DCAP8BWP7T $T=245160 413720 0 0 $X=244870 $Y=413485
X290 3 1 DCAP8BWP7T $T=248520 429400 1 0 $X=248230 $Y=425190
X291 3 1 DCAP8BWP7T $T=256360 476440 1 0 $X=256070 $Y=472230
X292 3 1 DCAP8BWP7T $T=274840 421560 1 0 $X=274550 $Y=417350
X293 3 1 DCAP8BWP7T $T=274840 429400 0 0 $X=274550 $Y=429165
X294 3 1 DCAP8BWP7T $T=276520 374520 0 0 $X=276230 $Y=374285
X295 3 1 DCAP8BWP7T $T=276520 390200 0 0 $X=276230 $Y=389965
X296 3 1 DCAP8BWP7T $T=282120 421560 1 0 $X=281830 $Y=417350
X297 3 1 DCAP8BWP7T $T=300040 413720 1 0 $X=299750 $Y=409510
X298 3 1 DCAP8BWP7T $T=301720 358840 0 0 $X=301430 $Y=358605
X299 3 1 DCAP8BWP7T $T=318520 358840 0 0 $X=318230 $Y=358605
X300 3 1 DCAP8BWP7T $T=318520 405880 1 0 $X=318230 $Y=401670
X301 3 1 DCAP8BWP7T $T=318520 413720 0 0 $X=318230 $Y=413485
X302 3 1 DCAP8BWP7T $T=318520 429400 1 0 $X=318230 $Y=425190
X303 3 1 DCAP8BWP7T $T=318520 429400 0 0 $X=318230 $Y=429165
X304 3 1 DCAP8BWP7T $T=318520 468600 0 0 $X=318230 $Y=468365
X305 3 1 DCAP8BWP7T $T=324120 382360 1 0 $X=323830 $Y=378150
X306 3 1 DCAP8BWP7T $T=347080 398040 0 0 $X=346790 $Y=397805
X307 3 1 DCAP8BWP7T $T=358840 476440 0 0 $X=358550 $Y=476205
X308 3 1 DCAP8BWP7T $T=360520 358840 0 0 $X=360230 $Y=358605
X309 3 1 DCAP8BWP7T $T=360520 366680 1 0 $X=360230 $Y=362470
X310 3 1 DCAP8BWP7T $T=360520 366680 0 0 $X=360230 $Y=366445
X311 3 1 DCAP8BWP7T $T=360520 382360 0 0 $X=360230 $Y=382125
X312 3 1 DCAP8BWP7T $T=360520 398040 1 0 $X=360230 $Y=393830
X313 3 1 DCAP8BWP7T $T=360520 421560 0 0 $X=360230 $Y=421325
X314 3 1 DCAP8BWP7T $T=360520 437240 1 0 $X=360230 $Y=433030
X315 3 1 DCAP8BWP7T $T=360520 437240 0 0 $X=360230 $Y=437005
X316 3 1 DCAP8BWP7T $T=360520 452920 1 0 $X=360230 $Y=448710
X317 3 1 DCAP8BWP7T $T=360520 460760 1 0 $X=360230 $Y=456550
X318 3 1 DCAP8BWP7T $T=366120 437240 0 0 $X=365830 $Y=437005
X319 3 1 DCAP8BWP7T $T=366120 468600 1 0 $X=365830 $Y=464390
X320 3 1 DCAP8BWP7T $T=366120 476440 0 0 $X=365830 $Y=476205
X321 3 1 DCAP8BWP7T $T=384040 382360 1 0 $X=383750 $Y=378150
X322 3 1 DCAP8BWP7T $T=386280 429400 0 0 $X=385990 $Y=429165
X323 3 1 DCAP8BWP7T $T=386840 413720 0 0 $X=386550 $Y=413485
X324 3 1 DCAP8BWP7T $T=390760 437240 0 0 $X=390470 $Y=437005
X325 3 1 DCAP8BWP7T $T=402520 437240 1 0 $X=402230 $Y=433030
X326 3 1 DCAP8BWP7T $T=402520 452920 1 0 $X=402230 $Y=448710
X327 3 1 DCAP8BWP7T $T=402520 460760 0 0 $X=402230 $Y=460525
X328 3 1 DCAP8BWP7T $T=402520 468600 0 0 $X=402230 $Y=468365
X329 3 1 DCAP8BWP7T $T=402520 484280 1 0 $X=402230 $Y=480070
X330 3 1 DCAP8BWP7T $T=412040 374520 0 0 $X=411750 $Y=374285
X331 3 1 DCAP8BWP7T $T=412600 413720 1 0 $X=412310 $Y=409510
X332 3 1 DCAP8BWP7T $T=426040 390200 1 0 $X=425750 $Y=385990
X333 3 1 DCAP8BWP7T $T=426040 476440 1 0 $X=425750 $Y=472230
X334 3 1 DCAP8BWP7T $T=428840 421560 0 0 $X=428550 $Y=421325
X335 3 1 DCAP8BWP7T $T=432760 398040 0 0 $X=432470 $Y=397805
X336 3 1 DCAP8BWP7T $T=442840 390200 1 0 $X=442550 $Y=385990
X337 3 1 DCAP8BWP7T $T=442840 460760 0 0 $X=442550 $Y=460525
X338 3 1 DCAP8BWP7T $T=443960 398040 1 0 $X=443670 $Y=393830
X339 3 1 DCAP8BWP7T $T=443960 413720 1 0 $X=443670 $Y=409510
X340 3 1 DCAP8BWP7T $T=443960 421560 0 0 $X=443670 $Y=421325
X341 3 1 DCAP8BWP7T $T=443960 468600 1 0 $X=443670 $Y=464390
X342 3 1 DCAP8BWP7T $T=444520 366680 1 0 $X=444230 $Y=362470
X343 3 1 DCAP8BWP7T $T=444520 398040 0 0 $X=444230 $Y=397805
X344 3 1 DCAP8BWP7T $T=444520 429400 1 0 $X=444230 $Y=425190
X345 3 1 DCAP8BWP7T $T=444520 437240 0 0 $X=444230 $Y=437005
X346 3 1 DCAP8BWP7T $T=444520 452920 0 0 $X=444230 $Y=452685
X347 3 1 DCAP8BWP7T $T=444520 468600 0 0 $X=444230 $Y=468365
X348 3 1 DCAP4BWP7T $T=156120 405880 0 0 $X=155830 $Y=405645
X349 3 1 DCAP4BWP7T $T=156120 445080 0 0 $X=155830 $Y=444845
X350 3 1 DCAP4BWP7T $T=156120 460760 1 0 $X=155830 $Y=456550
X351 3 1 DCAP4BWP7T $T=171800 476440 1 0 $X=171510 $Y=472230
X352 3 1 DCAP4BWP7T $T=172920 398040 1 0 $X=172630 $Y=393830
X353 3 1 DCAP4BWP7T $T=177400 437240 1 0 $X=177110 $Y=433030
X354 3 1 DCAP4BWP7T $T=183000 366680 0 0 $X=182710 $Y=366445
X355 3 1 DCAP4BWP7T $T=194200 398040 0 0 $X=193910 $Y=397805
X356 3 1 DCAP4BWP7T $T=194760 358840 0 0 $X=194470 $Y=358605
X357 3 1 DCAP4BWP7T $T=194760 398040 1 0 $X=194470 $Y=393830
X358 3 1 DCAP4BWP7T $T=194760 429400 0 0 $X=194470 $Y=429165
X359 3 1 DCAP4BWP7T $T=194760 476440 1 0 $X=194470 $Y=472230
X360 3 1 DCAP4BWP7T $T=207080 405880 1 0 $X=206790 $Y=401670
X361 3 1 DCAP4BWP7T $T=236200 374520 0 0 $X=235910 $Y=374285
X362 3 1 DCAP4BWP7T $T=236200 398040 0 0 $X=235910 $Y=397805
X363 3 1 DCAP4BWP7T $T=236760 358840 0 0 $X=236470 $Y=358605
X364 3 1 DCAP4BWP7T $T=236760 405880 1 0 $X=236470 $Y=401670
X365 3 1 DCAP4BWP7T $T=267000 445080 0 0 $X=266710 $Y=444845
X366 3 1 DCAP4BWP7T $T=278200 413720 0 0 $X=277910 $Y=413485
X367 3 1 DCAP4BWP7T $T=278200 421560 0 0 $X=277910 $Y=421325
X368 3 1 DCAP4BWP7T $T=278200 437240 1 0 $X=277910 $Y=433030
X369 3 1 DCAP4BWP7T $T=278200 437240 0 0 $X=277910 $Y=437005
X370 3 1 DCAP4BWP7T $T=278760 460760 0 0 $X=278470 $Y=460525
X371 3 1 DCAP4BWP7T $T=291080 476440 0 0 $X=290790 $Y=476205
X372 3 1 DCAP4BWP7T $T=299480 429400 1 0 $X=299190 $Y=425190
X373 3 1 DCAP4BWP7T $T=306760 390200 1 0 $X=306470 $Y=385990
X374 3 1 DCAP4BWP7T $T=320200 390200 0 0 $X=319910 $Y=389965
X375 3 1 DCAP4BWP7T $T=324120 382360 0 0 $X=323830 $Y=382125
X376 3 1 DCAP4BWP7T $T=324120 460760 0 0 $X=323830 $Y=460525
X377 3 1 DCAP4BWP7T $T=328600 437240 0 0 $X=328310 $Y=437005
X378 3 1 DCAP4BWP7T $T=331400 413720 1 0 $X=331110 $Y=409510
X379 3 1 DCAP4BWP7T $T=335320 460760 0 0 $X=335030 $Y=460525
X380 3 1 DCAP4BWP7T $T=345960 468600 1 0 $X=345670 $Y=464390
X381 3 1 DCAP4BWP7T $T=352120 476440 0 0 $X=351830 $Y=476205
X382 3 1 DCAP4BWP7T $T=362760 445080 1 0 $X=362470 $Y=440870
X383 3 1 DCAP4BWP7T $T=366120 358840 0 0 $X=365830 $Y=358605
X384 3 1 DCAP4BWP7T $T=366120 421560 0 0 $X=365830 $Y=421325
X385 3 1 DCAP4BWP7T $T=366120 429400 0 0 $X=365830 $Y=429165
X386 3 1 DCAP4BWP7T $T=379560 421560 0 0 $X=379270 $Y=421325
X387 3 1 DCAP4BWP7T $T=404200 429400 0 0 $X=403910 $Y=429165
X388 3 1 DCAP4BWP7T $T=404760 390200 1 0 $X=404470 $Y=385990
X389 3 1 DCAP4BWP7T $T=414280 421560 1 0 $X=413990 $Y=417350
X390 3 1 DCAP4BWP7T $T=423240 390200 0 0 $X=422950 $Y=389965
X391 3 1 ICV_40 $T=162840 405880 1 0 $X=162550 $Y=401670
X392 3 1 ICV_40 $T=162840 445080 1 0 $X=162550 $Y=440870
X393 3 1 ICV_40 $T=164520 484280 1 0 $X=164230 $Y=480070
X394 3 1 ICV_40 $T=165080 429400 1 0 $X=164790 $Y=425190
X395 3 1 ICV_40 $T=165080 437240 0 0 $X=164790 $Y=437005
X396 3 1 ICV_40 $T=171800 460760 0 0 $X=171510 $Y=460525
X397 3 1 ICV_40 $T=172920 421560 0 0 $X=172630 $Y=421325
X398 3 1 ICV_40 $T=188600 366680 1 0 $X=188310 $Y=362470
X399 3 1 ICV_40 $T=189720 460760 1 0 $X=189430 $Y=456550
X400 3 1 ICV_40 $T=190280 421560 0 0 $X=189990 $Y=421325
X401 3 1 ICV_40 $T=190280 452920 0 0 $X=189990 $Y=452685
X402 3 1 ICV_40 $T=207080 421560 0 0 $X=206790 $Y=421325
X403 3 1 ICV_40 $T=216040 460760 1 0 $X=215750 $Y=456550
X404 3 1 ICV_40 $T=230600 421560 0 0 $X=230310 $Y=421325
X405 3 1 ICV_40 $T=230600 460760 0 0 $X=230310 $Y=460525
X406 3 1 ICV_40 $T=231160 476440 0 0 $X=230870 $Y=476205
X407 3 1 ICV_40 $T=231720 382360 1 0 $X=231430 $Y=378150
X408 3 1 ICV_40 $T=231720 421560 1 0 $X=231430 $Y=417350
X409 3 1 ICV_40 $T=232280 366680 0 0 $X=231990 $Y=366445
X410 3 1 ICV_40 $T=242920 445080 1 0 $X=242630 $Y=440870
X411 3 1 ICV_40 $T=249080 429400 0 0 $X=248790 $Y=429165
X412 3 1 ICV_40 $T=272600 358840 0 0 $X=272310 $Y=358605
X413 3 1 ICV_40 $T=273720 484280 1 0 $X=273430 $Y=480070
X414 3 1 ICV_40 $T=274280 390200 1 0 $X=273990 $Y=385990
X415 3 1 ICV_40 $T=274280 398040 0 0 $X=273990 $Y=397805
X416 3 1 ICV_40 $T=282120 445080 0 0 $X=281830 $Y=444845
X417 3 1 ICV_40 $T=284360 382360 1 0 $X=284070 $Y=378150
X418 3 1 ICV_40 $T=286600 468600 0 0 $X=286310 $Y=468365
X419 3 1 ICV_40 $T=287720 374520 1 0 $X=287430 $Y=370310
X420 3 1 ICV_40 $T=294440 468600 1 0 $X=294150 $Y=464390
X421 3 1 ICV_40 $T=297240 398040 1 0 $X=296950 $Y=393830
X422 3 1 ICV_40 $T=315720 398040 1 0 $X=315430 $Y=393830
X423 3 1 ICV_40 $T=315720 398040 0 0 $X=315430 $Y=397805
X424 3 1 ICV_40 $T=315720 413720 1 0 $X=315430 $Y=409510
X425 3 1 ICV_40 $T=324120 476440 0 0 $X=323830 $Y=476205
X426 3 1 ICV_40 $T=349880 460760 1 0 $X=349590 $Y=456550
X427 3 1 ICV_40 $T=356600 468600 0 0 $X=356310 $Y=468365
X428 3 1 ICV_40 $T=357720 382360 1 0 $X=357430 $Y=378150
X429 3 1 ICV_40 $T=375080 452920 0 0 $X=374790 $Y=452685
X430 3 1 ICV_40 $T=378440 437240 0 0 $X=378150 $Y=437005
X431 3 1 ICV_40 $T=380680 468600 0 0 $X=380390 $Y=468365
X432 3 1 ICV_40 $T=390760 468600 0 0 $X=390470 $Y=468365
X433 3 1 ICV_40 $T=398600 421560 1 0 $X=398310 $Y=417350
X434 3 1 ICV_40 $T=399160 429400 1 0 $X=398870 $Y=425190
X435 3 1 ICV_40 $T=399720 476440 0 0 $X=399430 $Y=476205
X436 3 1 ICV_40 $T=400280 366680 0 0 $X=399990 $Y=366445
X437 3 1 ICV_40 $T=417080 437240 0 0 $X=416790 $Y=437005
X438 3 1 ICV_40 $T=417080 452920 1 0 $X=416790 $Y=448710
X439 3 1 ICV_40 $T=417080 452920 0 0 $X=416790 $Y=452685
X440 3 1 ICV_40 $T=426040 374520 1 0 $X=425750 $Y=370310
X441 3 1 ICV_40 $T=426040 413720 0 0 $X=425750 $Y=413485
X442 3 1 ICV_40 $T=433320 437240 0 0 $X=433030 $Y=437005
X443 3 1 ICV_40 $T=440600 405880 1 0 $X=440310 $Y=401670
X444 3 1 ICV_40 $T=441160 476440 0 0 $X=440870 $Y=476205
X445 3 1 ICV_40 $T=442280 382360 0 0 $X=441990 $Y=382125
X446 290 1 291 295 3 NR2D1BWP7T $T=156680 421560 1 0 $X=156390 $Y=417350
X447 297 1 303 299 3 NR2D1BWP7T $T=162280 460760 0 180 $X=159750 $Y=456550
X448 301 1 289 299 3 NR2D1BWP7T $T=160600 445080 1 0 $X=160310 $Y=440870
X449 290 1 305 302 3 NR2D1BWP7T $T=162840 445080 1 180 $X=160310 $Y=444845
X450 297 1 307 14 3 NR2D1BWP7T $T=160600 460760 0 0 $X=160310 $Y=460525
X451 295 1 308 14 3 NR2D1BWP7T $T=160600 468600 0 0 $X=160310 $Y=468365
X452 15 1 293 10 3 NR2D1BWP7T $T=163960 398040 0 180 $X=161430 $Y=393830
X453 290 1 313 301 3 NR2D1BWP7T $T=161720 421560 1 0 $X=161430 $Y=417350
X454 301 1 316 309 3 NR2D1BWP7T $T=162280 460760 1 0 $X=161990 $Y=456550
X455 301 1 315 14 3 NR2D1BWP7T $T=165080 445080 1 180 $X=162550 $Y=444845
X456 297 1 317 309 3 NR2D1BWP7T $T=162840 468600 0 0 $X=162550 $Y=468365
X457 301 1 319 304 3 NR2D1BWP7T $T=165080 421560 1 0 $X=164790 $Y=417350
X458 299 1 327 295 3 NR2D1BWP7T $T=169560 468600 0 0 $X=169270 $Y=468365
X459 311 1 320 14 3 NR2D1BWP7T $T=172920 421560 1 180 $X=170390 $Y=421325
X460 290 1 336 297 3 NR2D1BWP7T $T=175720 429400 0 180 $X=173190 $Y=425190
X461 311 1 338 290 3 NR2D1BWP7T $T=176840 429400 1 180 $X=174310 $Y=429165
X462 311 1 342 309 3 NR2D1BWP7T $T=177400 437240 0 180 $X=174870 $Y=433030
X463 311 1 344 299 3 NR2D1BWP7T $T=175720 421560 1 0 $X=175430 $Y=417350
X464 299 1 349 302 3 NR2D1BWP7T $T=176280 468600 0 0 $X=175990 $Y=468365
X465 398 1 400 73 3 NR2D1BWP7T $T=228360 421560 0 0 $X=228070 $Y=421325
X466 77 1 403 405 3 NR2D1BWP7T $T=230600 437240 1 0 $X=230310 $Y=433030
X467 405 1 425 97 3 NR2D1BWP7T $T=257480 437240 1 180 $X=254950 $Y=437005
X468 77 1 428 398 3 NR2D1BWP7T $T=257480 429400 1 0 $X=257190 $Y=425190
X469 429 1 446 73 3 NR2D1BWP7T $T=259720 405880 1 0 $X=259430 $Y=401670
X470 429 1 432 97 3 NR2D1BWP7T $T=261960 452920 0 180 $X=259430 $Y=448710
X471 77 1 435 429 3 NR2D1BWP7T $T=262520 413720 0 0 $X=262230 $Y=413485
X472 405 1 426 73 3 NR2D1BWP7T $T=265320 398040 1 180 $X=262790 $Y=397805
X473 405 1 442 105 3 NR2D1BWP7T $T=269240 366680 0 180 $X=266710 $Y=362470
X474 106 1 422 97 3 NR2D1BWP7T $T=269240 413720 1 180 $X=266710 $Y=413485
X475 398 1 430 97 3 NR2D1BWP7T $T=270360 421560 0 180 $X=267830 $Y=417350
X476 109 1 431 105 3 NR2D1BWP7T $T=271480 366680 0 180 $X=268950 $Y=362470
X477 109 1 452 110 3 NR2D1BWP7T $T=273720 366680 0 180 $X=271190 $Y=362470
X478 109 1 466 77 3 NR2D1BWP7T $T=287160 468600 0 180 $X=284630 $Y=464390
X479 119 1 123 122 3 NR2D1BWP7T $T=287720 374520 0 180 $X=285190 $Y=370310
X480 429 1 472 105 3 NR2D1BWP7T $T=291080 445080 1 180 $X=288550 $Y=444845
X481 429 1 476 131 3 NR2D1BWP7T $T=291080 429400 1 0 $X=290790 $Y=425190
X482 405 1 478 131 3 NR2D1BWP7T $T=294440 468600 0 180 $X=291910 $Y=464390
X483 105 1 483 398 3 NR2D1BWP7T $T=293320 429400 1 0 $X=293030 $Y=425190
X484 429 1 486 110 3 NR2D1BWP7T $T=295000 398040 1 0 $X=294710 $Y=393830
X485 398 1 487 110 3 NR2D1BWP7T $T=297240 429400 1 0 $X=296950 $Y=425190
X486 405 1 475 110 3 NR2D1BWP7T $T=304520 398040 1 0 $X=304230 $Y=393830
X487 109 1 489 131 3 NR2D1BWP7T $T=307880 468600 0 180 $X=305350 $Y=464390
X488 77 1 479 507 3 NR2D1BWP7T $T=307880 468600 0 0 $X=307590 $Y=468365
X489 109 1 495 514 3 NR2D1BWP7T $T=314600 468600 0 0 $X=314310 $Y=468365
X490 514 1 517 405 3 NR2D1BWP7T $T=318520 429400 0 180 $X=315990 $Y=425190
X491 105 1 506 507 3 NR2D1BWP7T $T=316280 429400 0 0 $X=315990 $Y=429165
X492 507 1 509 73 3 NR2D1BWP7T $T=326360 460760 0 0 $X=326070 $Y=460525
X493 150 1 151 10 3 NR2D1BWP7T $T=326920 413720 1 0 $X=326630 $Y=409510
X494 158 1 531 10 3 NR2D1BWP7T $T=329720 398040 0 180 $X=327190 $Y=393830
X495 77 1 484 540 3 NR2D1BWP7T $T=327480 460760 1 0 $X=327190 $Y=456550
X496 154 1 152 10 3 NR2D1BWP7T $T=330280 358840 1 180 $X=327750 $Y=358605
X497 507 1 155 97 3 NR2D1BWP7T $T=328040 468600 1 0 $X=327750 $Y=464390
X498 157 1 538 10 3 NR2D1BWP7T $T=331400 413720 0 180 $X=328870 $Y=409510
X499 540 1 159 97 3 NR2D1BWP7T $T=329720 460760 1 0 $X=329430 $Y=456550
X500 540 1 539 73 3 NR2D1BWP7T $T=335320 460760 1 180 $X=332790 $Y=460525
X501 162 1 546 163 3 NR2D1BWP7T $T=335880 390200 1 0 $X=335590 $Y=385990
X502 141 1 166 568 3 NR2D1BWP7T $T=340920 390200 1 0 $X=340630 $Y=385990
X503 568 1 566 10 3 NR2D1BWP7T $T=359400 374520 1 180 $X=356870 $Y=374285
X504 179 1 182 183 3 NR2D1BWP7T $T=358280 358840 0 0 $X=357990 $Y=358605
X505 180 1 561 569 3 NR2D1BWP7T $T=358280 460760 1 0 $X=357990 $Y=456550
X506 198 1 578 97 3 NR2D1BWP7T $T=374520 429400 1 180 $X=371990 $Y=429165
X507 183 1 565 10 3 NR2D1BWP7T $T=375640 398040 0 180 $X=373110 $Y=393830
X508 201 1 581 97 3 NR2D1BWP7T $T=375640 437240 1 180 $X=373110 $Y=437005
X509 588 1 580 97 3 NR2D1BWP7T $T=380680 437240 0 180 $X=378150 $Y=433030
X510 188 1 589 201 3 NR2D1BWP7T $T=385160 445080 0 180 $X=382630 $Y=440870
X511 174 1 590 97 3 NR2D1BWP7T $T=386280 429400 1 180 $X=383750 $Y=429165
X512 175 1 576 588 3 NR2D1BWP7T $T=386280 437240 0 0 $X=385990 $Y=437005
X513 174 1 593 209 3 NR2D1BWP7T $T=387960 445080 1 0 $X=387670 $Y=440870
X514 175 1 591 198 3 NR2D1BWP7T $T=390760 437240 1 180 $X=388230 $Y=437005
X515 209 1 599 201 3 NR2D1BWP7T $T=394680 445080 0 180 $X=392150 $Y=440870
X516 607 1 592 97 3 NR2D1BWP7T $T=396920 429400 0 180 $X=394390 $Y=425190
X517 609 1 214 97 3 NR2D1BWP7T $T=399160 429400 0 180 $X=396630 $Y=425190
X518 188 1 610 198 3 NR2D1BWP7T $T=400840 452920 0 180 $X=398310 $Y=448710
X519 174 1 601 220 3 NR2D1BWP7T $T=399160 452920 0 0 $X=398870 $Y=452685
X520 220 1 613 201 3 NR2D1BWP7T $T=401960 460760 0 180 $X=399430 $Y=456550
X521 175 1 617 609 3 NR2D1BWP7T $T=400280 437240 1 0 $X=399990 $Y=433030
X522 209 1 631 607 3 NR2D1BWP7T $T=408680 421560 0 0 $X=408390 $Y=421325
X523 188 1 606 588 3 NR2D1BWP7T $T=410920 445080 0 180 $X=408390 $Y=440870
X524 175 1 620 607 3 NR2D1BWP7T $T=409240 437240 1 0 $X=408950 $Y=433030
X525 209 1 626 588 3 NR2D1BWP7T $T=412040 445080 0 0 $X=411750 $Y=444845
X526 588 1 235 220 3 NR2D1BWP7T $T=416520 445080 1 180 $X=413990 $Y=444845
X527 220 1 619 198 3 NR2D1BWP7T $T=417640 445080 1 0 $X=417350 $Y=440870
X528 588 1 625 241 3 NR2D1BWP7T $T=418200 445080 0 0 $X=417910 $Y=444845
X529 188 1 636 607 3 NR2D1BWP7T $T=420440 437240 1 0 $X=420150 $Y=433030
X530 174 1 635 243 3 NR2D1BWP7T $T=426040 452920 0 180 $X=423510 $Y=448710
X531 243 1 644 201 3 NR2D1BWP7T $T=427720 452920 1 180 $X=425190 $Y=452685
X532 174 1 654 254 3 NR2D1BWP7T $T=430520 476440 1 0 $X=430230 $Y=472230
X533 609 1 652 188 3 NR2D1BWP7T $T=432760 445080 1 0 $X=432470 $Y=440870
X534 1 3 DCAP64BWP7T $T=198120 445080 1 0 $X=197830 $Y=440870
X535 1 3 DCAP64BWP7T $T=198120 468600 1 0 $X=197830 $Y=464390
X536 1 3 DCAP64BWP7T $T=198120 468600 0 0 $X=197830 $Y=468365
X537 1 3 DCAP64BWP7T $T=240120 398040 1 0 $X=239830 $Y=393830
X538 1 3 DCAP64BWP7T $T=240120 468600 0 0 $X=239830 $Y=468365
X539 1 3 DCAP64BWP7T $T=282120 366680 0 0 $X=281830 $Y=366445
X540 1 3 DCAP64BWP7T $T=282120 382360 0 0 $X=281830 $Y=382125
X541 1 3 DCAP64BWP7T $T=282120 421560 0 0 $X=281830 $Y=421325
X542 1 3 DCAP64BWP7T $T=282120 437240 1 0 $X=281830 $Y=433030
X543 1 3 DCAP64BWP7T $T=324120 476440 1 0 $X=323830 $Y=472230
X544 1 3 DCAP64BWP7T $T=328040 390200 0 0 $X=327750 $Y=389965
X545 1 3 DCAP64BWP7T $T=366120 405880 1 0 $X=365830 $Y=401670
X546 1 3 DCAP64BWP7T $T=366120 476440 1 0 $X=365830 $Y=472230
X577 1 3 DCAP32BWP7T $T=173480 405880 1 0 $X=173190 $Y=401670
X578 1 3 DCAP32BWP7T $T=174040 445080 1 0 $X=173750 $Y=440870
X579 1 3 DCAP32BWP7T $T=175720 429400 1 0 $X=175430 $Y=425190
X580 1 3 DCAP32BWP7T $T=175720 484280 1 0 $X=175430 $Y=480070
X581 1 3 DCAP32BWP7T $T=176280 398040 0 0 $X=175990 $Y=397805
X582 1 3 DCAP32BWP7T $T=176840 358840 0 0 $X=176550 $Y=358605
X583 1 3 DCAP32BWP7T $T=176840 429400 0 0 $X=176550 $Y=429165
X584 1 3 DCAP32BWP7T $T=198120 382360 1 0 $X=197830 $Y=378150
X585 1 3 DCAP32BWP7T $T=198120 460760 1 0 $X=197830 $Y=456550
X586 1 3 DCAP32BWP7T $T=206520 390200 1 0 $X=206230 $Y=385990
X587 1 3 DCAP32BWP7T $T=209320 398040 0 0 $X=209030 $Y=397805
X588 1 3 DCAP32BWP7T $T=211560 374520 1 0 $X=211270 $Y=370310
X589 1 3 DCAP32BWP7T $T=217160 382360 0 0 $X=216870 $Y=382125
X590 1 3 DCAP32BWP7T $T=218840 358840 0 0 $X=218550 $Y=358605
X591 1 3 DCAP32BWP7T $T=219400 413720 1 0 $X=219110 $Y=409510
X592 1 3 DCAP32BWP7T $T=240120 421560 1 0 $X=239830 $Y=417350
X593 1 3 DCAP32BWP7T $T=246840 484280 1 0 $X=246550 $Y=480070
X594 1 3 DCAP32BWP7T $T=251320 437240 1 0 $X=251030 $Y=433030
X595 1 3 DCAP32BWP7T $T=251880 460760 0 0 $X=251590 $Y=460525
X596 1 3 DCAP32BWP7T $T=263080 374520 1 0 $X=262790 $Y=370310
X597 1 3 DCAP32BWP7T $T=282120 460760 1 0 $X=281830 $Y=456550
X598 1 3 DCAP32BWP7T $T=289960 366680 1 0 $X=289670 $Y=362470
X599 1 3 DCAP32BWP7T $T=289960 421560 1 0 $X=289670 $Y=417350
X600 1 3 DCAP32BWP7T $T=294440 382360 1 0 $X=294150 $Y=378150
X601 1 3 DCAP32BWP7T $T=296120 429400 0 0 $X=295830 $Y=429165
X602 1 3 DCAP32BWP7T $T=326360 437240 1 0 $X=326070 $Y=433030
X603 1 3 DCAP32BWP7T $T=330840 366680 0 0 $X=330550 $Y=366445
X604 1 3 DCAP32BWP7T $T=331960 460760 1 0 $X=331670 $Y=456550
X605 1 3 DCAP32BWP7T $T=342600 366680 1 0 $X=342310 $Y=362470
X606 1 3 DCAP32BWP7T $T=366120 382360 1 0 $X=365830 $Y=378150
X607 1 3 DCAP32BWP7T $T=368920 413720 0 0 $X=368630 $Y=413485
X608 1 3 DCAP32BWP7T $T=380680 421560 1 0 $X=380390 $Y=417350
X609 1 3 DCAP32BWP7T $T=381240 405880 0 0 $X=380950 $Y=405645
X610 1 3 DCAP32BWP7T $T=387400 398040 1 0 $X=387110 $Y=393830
X611 1 3 DCAP32BWP7T $T=408120 366680 1 0 $X=407830 $Y=362470
X612 1 3 DCAP32BWP7T $T=408120 476440 1 0 $X=407830 $Y=472230
X613 1 3 DCAP32BWP7T $T=408120 476440 0 0 $X=407830 $Y=476205
X614 1 3 DCAP32BWP7T $T=421560 460760 1 0 $X=421270 $Y=456550
X615 1 3 DCAP32BWP7T $T=424360 382360 0 0 $X=424070 $Y=382125
X616 1 3 DCAP32BWP7T $T=427160 374520 0 0 $X=426870 $Y=374285
X617 1 3 DCAP32BWP7T $T=427720 484280 1 0 $X=427430 $Y=480070
X618 1 3 DCAP32BWP7T $T=429960 358840 0 0 $X=429670 $Y=358605
X619 1 3 DCAP32BWP7T $T=429960 452920 1 0 $X=429670 $Y=448710
X620 289 291 320 322 1 3 324 FA1D0BWP7T $T=156120 429400 0 0 $X=155830 $Y=429165
X621 17 316 32 347 1 3 35 FA1D0BWP7T $T=167880 460760 1 0 $X=167590 $Y=456550
X622 346 332 353 352 1 3 357 FA1D0BWP7T $T=178520 405880 0 0 $X=178230 $Y=405645
X623 305 303 342 356 1 3 355 FA1D0BWP7T $T=179080 445080 0 0 $X=178790 $Y=444845
X624 348 322 331 358 1 3 361 FA1D0BWP7T $T=179640 437240 1 0 $X=179350 $Y=433030
X625 308 349 317 359 1 3 45 FA1D0BWP7T $T=179640 460760 0 0 $X=179350 $Y=460525
X626 335 347 355 360 1 3 362 FA1D0BWP7T $T=179640 476440 0 0 $X=179350 $Y=476205
X627 300 319 336 363 1 3 375 FA1D0BWP7T $T=198680 421560 1 0 $X=198390 $Y=417350
X628 356 324 369 370 1 3 376 FA1D0BWP7T $T=198680 437240 1 0 $X=198390 $Y=433030
X629 329 326 315 369 1 3 385 FA1D0BWP7T $T=198680 452920 1 0 $X=198390 $Y=448710
X630 328 307 327 371 1 3 377 FA1D0BWP7T $T=198680 460760 0 0 $X=198390 $Y=460525
X631 46 365 362 372 1 3 62 FA1D0BWP7T $T=198680 476440 0 0 $X=198390 $Y=476205
X632 360 371 385 389 1 3 381 FA1D0BWP7T $T=207080 445080 0 0 $X=206790 $Y=444845
X633 54 57 384 65 1 3 374 FA1D0BWP7T $T=210440 366680 0 0 $X=210150 $Y=366445
X634 394 372 381 380 1 3 378 FA1D0BWP7T $T=224440 437240 0 180 $X=211270 $Y=433030
X635 359 377 58 365 1 3 379 FA1D0BWP7T $T=224440 460760 1 180 $X=211270 $Y=460525
X636 67 395 79 80 1 3 82 FA1D0BWP7T $T=221640 366680 1 0 $X=221350 $Y=362470
X637 361 393 370 406 1 3 407 FA1D0BWP7T $T=221640 405880 0 0 $X=221350 $Y=405645
X638 423 426 435 441 1 3 445 FA1D0BWP7T $T=252440 390200 1 0 $X=252150 $Y=385990
X639 433 448 444 456 1 3 401 FA1D0BWP7T $T=263640 374520 0 0 $X=263350 $Y=374285
X640 442 428 452 457 1 3 459 FA1D0BWP7T $T=263640 390200 0 0 $X=263350 $Y=389965
X641 462 457 453 463 1 3 460 FA1D0BWP7T $T=295560 390200 1 180 $X=282390 $Y=389965
X642 451 465 475 481 1 3 485 FA1D0BWP7T $T=282680 405880 1 0 $X=282390 $Y=401670
X643 464 486 483 493 1 3 497 FA1D0BWP7T $T=292760 413720 0 0 $X=292470 $Y=413485
X644 479 472 489 482 1 3 498 FA1D0BWP7T $T=292760 445080 1 0 $X=292470 $Y=440870
X645 460 480 494 496 1 3 502 FA1D0BWP7T $T=293880 390200 1 0 $X=293590 $Y=385990
X646 482 459 481 494 1 3 503 FA1D0BWP7T $T=293880 398040 0 0 $X=293590 $Y=397805
X647 484 478 495 504 1 3 501 FA1D0BWP7T $T=295000 452920 0 0 $X=294710 $Y=452685
X648 487 506 476 490 1 3 488 FA1D0BWP7T $T=314600 429400 0 180 $X=301430 $Y=425190
X649 500 493 485 515 1 3 520 FA1D0BWP7T $T=305640 405880 1 0 $X=305350 $Y=401670
X650 490 497 512 516 1 3 521 FA1D0BWP7T $T=305640 413720 0 0 $X=305350 $Y=413485
X651 499 504 498 500 1 3 522 FA1D0BWP7T $T=305640 445080 1 0 $X=305350 $Y=440870
X652 501 505 513 518 1 3 523 FA1D0BWP7T $T=305640 460760 1 0 $X=305350 $Y=456550
X653 541 548 520 543 1 3 547 FA1D0BWP7T $T=334200 398040 0 0 $X=333910 $Y=397805
X654 518 516 522 548 1 3 533 FA1D0BWP7T $T=350440 429400 0 180 $X=337270 $Y=425190
X655 517 562 532 512 1 3 544 FA1D0BWP7T $T=360520 421560 1 180 $X=347350 $Y=421325
X656 574 579 585 195 1 3 206 FA1D0BWP7T $T=369480 452920 1 0 $X=369190 $Y=448710
X657 577 582 586 569 1 3 189 FA1D0BWP7T $T=371160 468600 1 0 $X=370870 $Y=464390
X658 570 589 593 595 1 3 200 FA1D0BWP7T $T=377880 476440 0 0 $X=377590 $Y=476205
X659 606 601 591 579 1 3 208 FA1D0BWP7T $T=395240 452920 1 180 $X=382070 $Y=452685
X660 598 604 610 221 1 3 224 FA1D0BWP7T $T=389640 484280 1 0 $X=389350 $Y=480070
X661 619 625 631 239 1 3 242 FA1D0BWP7T $T=408680 460760 1 0 $X=408390 $Y=456550
X662 240 626 620 229 1 3 226 FA1D0BWP7T $T=421560 468600 1 180 $X=408390 $Y=468365
X663 635 636 617 255 1 3 257 FA1D0BWP7T $T=421000 460760 0 0 $X=420710 $Y=460525
X664 652 654 659 273 1 3 278 FA1D0BWP7T $T=431640 468600 0 0 $X=431350 $Y=468365
X665 292 3 1 297 INVD1BWP7T $T=158360 460760 1 0 $X=158070 $Y=456550
X666 11 3 1 304 INVD1BWP7T $T=161160 476440 1 0 $X=160870 $Y=472230
X667 12 3 1 311 INVD1BWP7T $T=170680 421560 1 0 $X=170390 $Y=417350
X668 21 3 1 299 INVD1BWP7T $T=171240 484280 1 0 $X=170950 $Y=480070
X669 24 3 1 290 INVD1BWP7T $T=173480 445080 1 180 $X=171510 $Y=444845
X670 23 3 1 301 INVD1BWP7T $T=173480 437240 0 0 $X=173190 $Y=437005
X671 38 3 1 39 INVD1BWP7T $T=185240 366680 0 0 $X=184950 $Y=366445
X672 74 3 1 325 INVD1BWP7T $T=230600 437240 0 180 $X=228630 $Y=433030
X673 455 3 1 429 INVD1BWP7T $T=290520 413720 1 180 $X=288550 $Y=413485
X674 470 3 1 105 INVD1BWP7T $T=296120 429400 1 180 $X=294150 $Y=429165
X675 471 3 1 398 INVD1BWP7T $T=297240 429400 0 180 $X=295270 $Y=425190
X676 144 3 1 131 INVD1BWP7T $T=318520 468600 1 180 $X=316550 $Y=468365
X677 527 3 1 110 INVD1BWP7T $T=326360 437240 0 180 $X=324390 $Y=433030
X678 530 3 1 514 INVD1BWP7T $T=328600 452920 0 180 $X=326630 $Y=448710
X679 529 3 1 507 INVD1BWP7T $T=334200 476440 1 180 $X=332230 $Y=476205
X680 213 3 1 607 INVD1BWP7T $T=397480 413720 0 180 $X=395510 $Y=409510
X681 203 3 1 588 INVD1BWP7T $T=399160 445080 0 180 $X=397190 $Y=440870
X682 207 3 1 201 INVD1BWP7T $T=399720 468600 1 0 $X=399430 $Y=464390
X683 223 3 1 220 INVD1BWP7T $T=402520 452920 0 180 $X=400550 $Y=448710
X684 211 3 1 209 INVD1BWP7T $T=414280 445080 0 180 $X=412310 $Y=440870
X685 643 3 1 243 INVD1BWP7T $T=426040 468600 0 0 $X=425750 $Y=468365
X686 629 3 1 241 INVD1BWP7T $T=429400 421560 1 0 $X=429110 $Y=417350
X801 292 3 296 11 1 ND2D1BWP7T $T=158360 405880 0 0 $X=158070 $Y=405645
X802 12 3 306 11 1 ND2D1BWP7T $T=160600 405880 1 0 $X=160310 $Y=401670
X803 7 3 318 11 1 ND2D1BWP7T $T=161160 452920 0 0 $X=160870 $Y=452685
X804 292 3 314 16 1 ND2D1BWP7T $T=162280 484280 1 0 $X=161990 $Y=480070
X805 27 3 339 26 1 ND2D1BWP7T $T=174600 358840 0 0 $X=174310 $Y=358605
X806 30 3 343 33 1 ND2D1BWP7T $T=175160 398040 1 0 $X=174870 $Y=393830
X807 48 3 364 31 1 ND2D1BWP7T $T=202600 405880 1 180 $X=200070 $Y=405645
X808 59 3 373 60 1 ND2D1BWP7T $T=216600 358840 0 0 $X=216310 $Y=358605
X809 411 3 399 24 1 ND2D1BWP7T $T=242920 445080 0 180 $X=240390 $Y=440870
X810 96 3 420 69 1 ND2D1BWP7T $T=254680 374520 1 180 $X=252150 $Y=374285
X811 114 3 438 112 1 ND2D1BWP7T $T=275400 452920 0 180 $X=272870 $Y=448710
X812 138 3 526 458 1 ND2D1BWP7T $T=324680 413720 1 0 $X=324390 $Y=409510
X813 471 3 524 144 1 ND2D1BWP7T $T=324680 445080 1 0 $X=324390 $Y=440870
X814 470 3 534 535 1 ND2D1BWP7T $T=327480 445080 0 0 $X=327190 $Y=444845
X815 146 3 525 156 1 ND2D1BWP7T $T=328600 382360 1 0 $X=328310 $Y=378150
X816 563 3 553 454 1 ND2D1BWP7T $T=354360 445080 1 180 $X=351830 $Y=444845
X817 559 3 550 112 1 ND2D1BWP7T $T=353240 452920 1 0 $X=352950 $Y=448710
X818 529 3 554 527 1 ND2D1BWP7T $T=360520 437240 0 180 $X=357990 $Y=433030
X819 455 3 564 530 1 ND2D1BWP7T $T=368920 413720 1 180 $X=366390 $Y=413485
X820 193 3 556 114 1 ND2D1BWP7T $T=379000 413720 0 180 $X=376470 $Y=409510
X821 202 3 575 207 1 ND2D1BWP7T $T=380680 445080 1 0 $X=380390 $Y=440870
X822 202 3 247 217 1 ND2D1BWP7T $T=424920 437240 0 0 $X=424630 $Y=437005
X823 262 3 647 261 1 ND2D1BWP7T $T=439480 445080 0 180 $X=436950 $Y=440870
X842 9 3 1 302 INVD0BWP7T $T=159480 476440 1 0 $X=159190 $Y=472230
X843 13 3 1 309 INVD0BWP7T $T=160600 484280 1 0 $X=160310 $Y=480070
X844 52 3 1 333 INVD0BWP7T $T=176840 437240 1 180 $X=174870 $Y=437005
X845 334 3 1 348 INVD0BWP7T $T=179640 421560 0 0 $X=179350 $Y=421325
X846 363 3 1 353 INVD0BWP7T $T=200360 405880 1 180 $X=198390 $Y=405645
X847 387 3 1 341 INVD0BWP7T $T=217720 421560 0 180 $X=215750 $Y=417350
X848 386 3 1 393 INVD0BWP7T $T=225000 390200 1 180 $X=223030 $Y=389965
X849 357 3 1 391 INVD0BWP7T $T=228920 429400 0 180 $X=226950 $Y=425190
X850 70 3 1 337 INVD0BWP7T $T=229480 476440 1 180 $X=227510 $Y=476205
X851 402 3 1 72 INVD0BWP7T $T=231160 476440 1 180 $X=229190 $Y=476205
X852 401 3 1 404 INVD0BWP7T $T=230040 374520 0 0 $X=229750 $Y=374285
X853 64 3 1 312 INVD0BWP7T $T=232840 390200 1 180 $X=230870 $Y=389965
X854 441 3 1 444 INVD0BWP7T $T=263640 366680 1 0 $X=263350 $Y=362470
X855 108 3 1 443 INVD0BWP7T $T=269240 476440 1 0 $X=268950 $Y=472230
X856 437 3 1 462 INVD0BWP7T $T=282680 382360 1 0 $X=282390 $Y=378150
X857 469 3 1 436 INVD0BWP7T $T=287720 452920 0 180 $X=285750 $Y=448710
X858 477 3 1 480 INVD0BWP7T $T=292760 382360 1 0 $X=292470 $Y=378150
X859 491 3 1 508 INVD0BWP7T $T=309560 390200 0 0 $X=309270 $Y=389965
X860 535 3 1 540 INVD0BWP7T $T=339240 460760 1 180 $X=337270 $Y=460525
X861 571 3 1 574 INVD0BWP7T $T=366680 445080 1 0 $X=366390 $Y=440870
X862 195 3 1 196 INVD0BWP7T $T=370600 476440 0 0 $X=370310 $Y=476205
X863 200 3 1 194 INVD0BWP7T $T=373960 476440 1 180 $X=371990 $Y=476205
X864 595 3 1 586 INVD0BWP7T $T=390760 468600 1 180 $X=388790 $Y=468365
X865 216 3 1 568 INVD0BWP7T $T=400280 366680 1 180 $X=398310 $Y=366445
X866 260 3 1 609 INVD0BWP7T $T=437240 445080 0 180 $X=435270 $Y=440870
X867 344 346 34 334 3 1 OAI21D0BWP7T $T=177960 421560 1 0 $X=177670 $Y=417350
X868 95 424 98 99 3 1 OAI21D0BWP7T $T=253560 476440 1 0 $X=253270 $Y=472230
X869 376 416 389 407 3 1 OAI21D0BWP7T $T=254680 429400 1 0 $X=254390 $Y=425190
X870 431 433 434 437 3 1 OAI21D0BWP7T $T=260280 374520 1 0 $X=259990 $Y=370310
X871 503 528 515 502 3 1 OAI21D0BWP7T $T=328040 398040 1 180 $X=324950 $Y=397805
X872 576 577 181 571 3 1 OAI21D0BWP7T $T=370600 437240 0 0 $X=370310 $Y=437005
X873 233 587 218 612 3 1 OAI21D0BWP7T $T=402520 382360 1 180 $X=399430 $Y=382125
X874 218 600 227 622 3 1 OAI21D0BWP7T $T=408680 390200 0 0 $X=408390 $Y=389965
X875 232 605 227 616 3 1 OAI21D0BWP7T $T=411480 405880 1 180 $X=408390 $Y=405645
X876 228 621 232 623 3 1 OAI21D0BWP7T $T=409800 413720 1 0 $X=409510 $Y=409510
X877 230 603 232 624 3 1 OAI21D0BWP7T $T=410360 366680 0 0 $X=410070 $Y=366445
X878 233 602 232 627 3 1 OAI21D0BWP7T $T=411480 382360 0 0 $X=411190 $Y=382125
X879 228 632 218 628 3 1 OAI21D0BWP7T $T=418760 398040 1 180 $X=415670 $Y=397805
X880 228 641 245 645 3 1 OAI21D0BWP7T $T=423240 413720 1 0 $X=422950 $Y=409510
X881 243 650 588 647 3 1 OAI21D0BWP7T $T=425480 445080 0 0 $X=425190 $Y=444845
X882 245 649 227 638 3 1 OAI21D0BWP7T $T=432760 398040 1 180 $X=429670 $Y=397805
X883 230 640 245 642 3 1 OAI21D0BWP7T $T=436120 374520 0 180 $X=433030 $Y=370310
X884 233 653 245 639 3 1 OAI21D0BWP7T $T=436120 390200 0 180 $X=433030 $Y=385990
X885 250 646 245 651 3 1 OAI21D0BWP7T $T=438920 366680 1 180 $X=435830 $Y=366445
X886 274 655 227 656 3 1 OAI21D0BWP7T $T=444520 398040 1 180 $X=441430 $Y=397805
X887 228 658 274 279 3 1 OAI21D0BWP7T $T=441720 413720 0 0 $X=441430 $Y=413485
X888 241 271 198 277 3 1 OAI21D0BWP7T $T=441720 429400 1 0 $X=441430 $Y=425190
X925 26 3 28 31 1 340 ND3D0BWP7T $T=173480 398040 0 0 $X=173190 $Y=397805
X926 34 3 12 21 1 334 ND3D0BWP7T $T=176280 445080 1 180 $X=173190 $Y=444845
X927 75 3 12 24 1 387 ND3D0BWP7T $T=230600 460760 1 180 $X=227510 $Y=460525
X928 434 3 114 470 1 437 ND3D0BWP7T $T=286040 413720 0 0 $X=285750 $Y=413485
X929 117 3 114 454 1 469 ND3D0BWP7T $T=290520 452920 0 180 $X=287430 $Y=448710
X930 153 3 535 112 1 542 ND3D0BWP7T $T=360520 452920 0 180 $X=357430 $Y=448710
X931 181 3 202 203 1 571 ND3D0BWP7T $T=375640 437240 0 0 $X=375350 $Y=437005
X932 251 3 643 207 1 249 ND3D0BWP7T $T=429400 476440 0 0 $X=429110 $Y=476205
X933 3 1 DCAP16BWP7T $T=163960 398040 1 0 $X=163670 $Y=393830
X934 3 1 DCAP16BWP7T $T=163960 413720 0 0 $X=163670 $Y=413485
X935 3 1 DCAP16BWP7T $T=174040 366680 0 0 $X=173750 $Y=366445
X936 3 1 DCAP16BWP7T $T=177400 398040 1 0 $X=177110 $Y=393830
X937 3 1 DCAP16BWP7T $T=179640 366680 1 0 $X=179350 $Y=362470
X938 3 1 DCAP16BWP7T $T=180760 460760 1 0 $X=180470 $Y=456550
X939 3 1 DCAP16BWP7T $T=181320 452920 0 0 $X=181030 $Y=452685
X940 3 1 DCAP16BWP7T $T=198120 413720 1 0 $X=197830 $Y=409510
X941 3 1 DCAP16BWP7T $T=216040 374520 0 0 $X=215750 $Y=374285
X942 3 1 DCAP16BWP7T $T=216040 429400 0 0 $X=215750 $Y=429165
X943 3 1 DCAP16BWP7T $T=218280 421560 0 0 $X=217990 $Y=421325
X944 3 1 DCAP16BWP7T $T=223320 366680 0 0 $X=223030 $Y=366445
X945 3 1 DCAP16BWP7T $T=227240 398040 0 0 $X=226950 $Y=397805
X946 3 1 DCAP16BWP7T $T=228920 429400 1 0 $X=228630 $Y=425190
X947 3 1 DCAP16BWP7T $T=229480 374520 1 0 $X=229190 $Y=370310
X948 3 1 DCAP16BWP7T $T=229480 452920 1 0 $X=229190 $Y=448710
X949 3 1 DCAP16BWP7T $T=240120 452920 0 0 $X=239830 $Y=452685
X950 3 1 DCAP16BWP7T $T=240120 468600 1 0 $X=239830 $Y=464390
X951 3 1 DCAP16BWP7T $T=251320 390200 0 0 $X=251030 $Y=389965
X952 3 1 DCAP16BWP7T $T=253560 366680 1 0 $X=253270 $Y=362470
X953 3 1 DCAP16BWP7T $T=258040 445080 0 0 $X=257750 $Y=444845
X954 3 1 DCAP16BWP7T $T=259720 429400 0 0 $X=259430 $Y=429165
X955 3 1 DCAP16BWP7T $T=261960 445080 1 0 $X=261670 $Y=440870
X956 3 1 DCAP16BWP7T $T=263640 358840 0 0 $X=263350 $Y=358605
X957 3 1 DCAP16BWP7T $T=264760 484280 1 0 $X=264470 $Y=480070
X958 3 1 DCAP16BWP7T $T=265320 390200 1 0 $X=265030 $Y=385990
X959 3 1 DCAP16BWP7T $T=265320 398040 0 0 $X=265030 $Y=397805
X960 3 1 DCAP16BWP7T $T=269240 413720 0 0 $X=268950 $Y=413485
X961 3 1 DCAP16BWP7T $T=269240 421560 0 0 $X=268950 $Y=421325
X962 3 1 DCAP16BWP7T $T=269240 437240 1 0 $X=268950 $Y=433030
X963 3 1 DCAP16BWP7T $T=269240 437240 0 0 $X=268950 $Y=437005
X964 3 1 DCAP16BWP7T $T=269800 460760 0 0 $X=269510 $Y=460525
X965 3 1 DCAP16BWP7T $T=271480 445080 0 0 $X=271190 $Y=444845
X966 3 1 DCAP16BWP7T $T=282120 398040 1 0 $X=281830 $Y=393830
X967 3 1 DCAP16BWP7T $T=282120 445080 1 0 $X=281830 $Y=440870
X968 3 1 DCAP16BWP7T $T=287160 484280 1 0 $X=286870 $Y=480070
X969 3 1 DCAP16BWP7T $T=293880 374520 0 0 $X=293590 $Y=374285
X970 3 1 DCAP16BWP7T $T=304520 484280 1 0 $X=304230 $Y=480070
X971 3 1 DCAP16BWP7T $T=306760 398040 1 0 $X=306470 $Y=393830
X972 3 1 DCAP16BWP7T $T=306760 398040 0 0 $X=306470 $Y=397805
X973 3 1 DCAP16BWP7T $T=310120 437240 0 0 $X=309830 $Y=437005
X974 3 1 DCAP16BWP7T $T=311240 390200 0 0 $X=310950 $Y=389965
X975 3 1 DCAP16BWP7T $T=312360 382360 1 0 $X=312070 $Y=378150
X976 3 1 DCAP16BWP7T $T=313480 374520 1 0 $X=313190 $Y=370310
X977 3 1 DCAP16BWP7T $T=324120 374520 1 0 $X=323830 $Y=370310
X978 3 1 DCAP16BWP7T $T=328600 382360 0 0 $X=328310 $Y=382125
X979 3 1 DCAP16BWP7T $T=339240 460760 0 0 $X=338950 $Y=460525
X980 3 1 DCAP16BWP7T $T=342040 452920 0 0 $X=341750 $Y=452685
X981 3 1 DCAP16BWP7T $T=346520 358840 0 0 $X=346230 $Y=358605
X982 3 1 DCAP16BWP7T $T=347640 468600 0 0 $X=347350 $Y=468365
X983 3 1 DCAP16BWP7T $T=348760 382360 1 0 $X=348470 $Y=378150
X984 3 1 DCAP16BWP7T $T=352120 460760 0 0 $X=351830 $Y=460525
X985 3 1 DCAP16BWP7T $T=354360 398040 0 0 $X=354070 $Y=397805
X986 3 1 DCAP16BWP7T $T=354360 445080 0 0 $X=354070 $Y=444845
X987 3 1 DCAP16BWP7T $T=354360 452920 0 0 $X=354070 $Y=452685
X988 3 1 DCAP16BWP7T $T=370600 421560 0 0 $X=370310 $Y=421325
X989 3 1 DCAP16BWP7T $T=371720 468600 0 0 $X=371430 $Y=468365
X990 3 1 DCAP16BWP7T $T=374520 429400 0 0 $X=374230 $Y=429165
X991 3 1 DCAP16BWP7T $T=379000 358840 0 0 $X=378710 $Y=358605
X992 3 1 DCAP16BWP7T $T=382920 429400 1 0 $X=382630 $Y=425190
X993 3 1 DCAP16BWP7T $T=389080 366680 0 0 $X=388790 $Y=366445
X994 3 1 DCAP16BWP7T $T=389080 382360 0 0 $X=388790 $Y=382125
X995 3 1 DCAP16BWP7T $T=389080 460760 0 0 $X=388790 $Y=460525
X996 3 1 DCAP16BWP7T $T=390760 476440 0 0 $X=390470 $Y=476205
X997 3 1 DCAP16BWP7T $T=397480 413720 1 0 $X=397190 $Y=409510
X998 3 1 DCAP16BWP7T $T=398040 437240 0 0 $X=397750 $Y=437005
X999 3 1 DCAP16BWP7T $T=411480 437240 1 0 $X=411190 $Y=433030
X1000 3 1 DCAP16BWP7T $T=419880 445080 1 0 $X=419590 $Y=440870
X1001 3 1 DCAP16BWP7T $T=431640 405880 1 0 $X=431350 $Y=401670
X1002 3 1 DCAP16BWP7T $T=436120 390200 0 0 $X=435830 $Y=389965
X1003 3 1 DCAP16BWP7T $T=438920 366680 0 0 $X=438630 $Y=366445
X1004 3 1 DCAP16BWP7T $T=438920 429400 0 0 $X=438630 $Y=429165
X1005 3 1 DCAP16BWP7T $T=439480 460760 1 0 $X=439190 $Y=456550
X1062 304 3 311 312 300 1 NR3D1BWP7T $T=159480 413720 0 0 $X=159190 $Y=413485
X1063 304 3 295 325 328 1 NR3D1BWP7T $T=171800 468600 0 0 $X=171510 $Y=468365
X1064 73 3 109 443 423 1 NR3D1BWP7T $T=275960 445080 0 180 $X=271190 $Y=440870
X1065 141 3 139 508 140 1 NR3D1BWP7T $T=310680 366680 1 0 $X=310390 $Y=362470
X1066 174 3 175 177 173 1 NR3D1BWP7T $T=358840 476440 1 180 $X=354070 $Y=476205
X1067 201 3 175 192 570 1 NR3D1BWP7T $T=384600 468600 1 0 $X=384310 $Y=464390
X1068 341 313 3 1 323 332 MAOI222D1BWP7T $T=175160 405880 1 180 $X=170390 $Y=405645
X1069 391 358 3 1 375 386 MAOI222D1BWP7T $T=218280 421560 1 180 $X=213510 $Y=421325
X1070 130 127 3 1 126 402 MAOI222D1BWP7T $T=291080 476440 1 180 $X=286310 $Y=476205
X1071 404 463 3 1 445 477 MAOI222D1BWP7T $T=309000 374520 1 0 $X=308710 $Y=370310
X1072 173 185 3 1 190 582 MAOI222D1BWP7T $T=366680 460760 0 0 $X=366390 $Y=460525
X1073 306 312 3 300 323 1 AOI21D1BWP7T $T=167320 405880 0 0 $X=167030 $Y=405645
X1074 325 318 3 328 326 1 AOI21D1BWP7T $T=168440 445080 0 0 $X=168150 $Y=444845
X1075 443 438 3 423 439 1 AOI21D1BWP7T $T=264760 437240 1 180 $X=261110 $Y=437005
X1076 454 77 1 3 INVD2BWP7T $T=271480 445080 1 180 $X=268950 $Y=444845
X1077 114 109 1 3 INVD2BWP7T $T=274840 405880 0 180 $X=272310 $Y=401670
X1078 112 73 1 3 INVD2BWP7T $T=274840 421560 0 180 $X=272310 $Y=417350
X1079 138 405 1 3 INVD2BWP7T $T=306760 413720 0 180 $X=304230 $Y=409510
X1080 146 139 1 3 INVD2BWP7T $T=325800 390200 0 0 $X=325510 $Y=389965
X1081 572 186 1 3 INVD2BWP7T $T=369480 405880 1 180 $X=366950 $Y=405645
X1082 202 175 1 3 INVD2BWP7T $T=395800 437240 0 0 $X=395510 $Y=437005
X1083 217 174 1 3 INVD2BWP7T $T=400280 460760 0 0 $X=399990 $Y=460525
X1148 5 8 3 1 321 DFQD0BWP7T $T=156680 366680 1 0 $X=156390 $Y=362470
X1149 5 6 3 1 294 DFQD0BWP7T $T=156680 374520 0 0 $X=156390 $Y=374285
X1150 5 19 3 1 298 DFQD0BWP7T $T=169000 366680 1 0 $X=168710 $Y=362470
X1151 5 20 3 1 330 DFQD0BWP7T $T=169000 374520 0 0 $X=168710 $Y=374285
X1152 5 36 3 1 33 DFQD0BWP7T $T=180760 374520 0 0 $X=180470 $Y=374285
X1153 61 396 3 1 81 DFQD0BWP7T $T=223880 476440 1 0 $X=223590 $Y=472230
X1154 5 418 3 1 60 DFQD0BWP7T $T=251320 390200 1 180 $X=240390 $Y=389965
X1155 5 413 3 1 92 DFQD0BWP7T $T=240680 405880 0 0 $X=240390 $Y=405645
X1156 61 419 3 1 84 DFQD0BWP7T $T=251320 437240 0 180 $X=240390 $Y=433030
X1157 61 427 3 1 411 DFQD0BWP7T $T=261960 445080 0 180 $X=251030 $Y=440870
X1158 5 103 3 1 408 DFQD0BWP7T $T=263640 358840 1 180 $X=252710 $Y=358605
X1159 61 425 3 1 440 DFQD0BWP7T $T=253000 452920 0 0 $X=252710 $Y=452685
X1160 61 447 3 1 108 DFQD0BWP7T $T=265320 452920 0 0 $X=265030 $Y=452685
X1161 61 432 3 1 417 DFQD0BWP7T $T=275960 468600 0 180 $X=265030 $Y=464390
X1162 61 473 3 1 117 DFQD0BWP7T $T=293320 452920 1 180 $X=282390 $Y=452685
X1163 142 510 3 1 137 DFQD0BWP7T $T=317960 374520 1 180 $X=307030 $Y=374285
X1164 142 511 3 1 491 DFQD0BWP7T $T=318520 358840 1 180 $X=307590 $Y=358605
X1165 61 537 3 1 492 DFQD0BWP7T $T=335320 484280 0 180 $X=324390 $Y=480070
X1166 61 168 3 1 530 DFQD0BWP7T $T=347640 468600 1 180 $X=336710 $Y=468365
X1167 61 167 3 1 527 DFQD0BWP7T $T=347640 484280 0 180 $X=336710 $Y=480070
X1168 142 545 3 1 552 DFQD0BWP7T $T=349880 382360 1 180 $X=338950 $Y=382125
X1169 61 561 3 1 181 DFQD0BWP7T $T=348760 484280 1 0 $X=348470 $Y=480070
X1170 142 565 3 1 558 DFQD0BWP7T $T=360520 366680 1 180 $X=349590 $Y=366445
X1171 142 567 3 1 557 DFQD0BWP7T $T=360520 398040 0 180 $X=349590 $Y=393830
X1172 142 580 3 1 184 DFQD0BWP7T $T=377320 374520 0 180 $X=366390 $Y=370310
X1173 142 578 3 1 572 DFQD0BWP7T $T=381240 405880 1 180 $X=370310 $Y=405645
X1174 142 590 3 1 583 DFQD0BWP7T $T=387400 398040 0 180 $X=376470 $Y=393830
X1175 142 592 3 1 204 DFQD0BWP7T $T=389080 366680 1 180 $X=378150 $Y=366445
X1176 142 587 3 1 594 DFQD0BWP7T $T=378440 382360 0 0 $X=378150 $Y=382125
X1177 142 596 3 1 205 DFQD0BWP7T $T=392440 413720 0 180 $X=381510 $Y=409510
X1178 142 597 3 1 573 DFQD0BWP7T $T=392440 421560 1 180 $X=381510 $Y=421325
X1179 142 600 3 1 608 DFQD0BWP7T $T=387960 398040 0 0 $X=387670 $Y=397805
X1180 142 602 3 1 611 DFQD0BWP7T $T=389640 390200 1 0 $X=389350 $Y=385990
X1181 142 603 3 1 615 DFQD0BWP7T $T=390760 374520 1 0 $X=390470 $Y=370310
X1182 142 210 3 1 618 DFQD0BWP7T $T=391880 358840 0 0 $X=391590 $Y=358605
X1183 142 605 3 1 614 DFQD0BWP7T $T=391880 413720 0 0 $X=391590 $Y=413485
X1184 142 640 3 1 630 DFQD0BWP7T $T=427160 374520 1 180 $X=416230 $Y=374285
X1185 142 632 3 1 629 DFQD0BWP7T $T=416520 421560 1 0 $X=416230 $Y=417350
X1186 142 646 3 1 633 DFQD0BWP7T $T=429960 358840 1 180 $X=419030 $Y=358605
X1187 142 649 3 1 634 DFQD0BWP7T $T=431640 405880 0 180 $X=420710 $Y=401670
X1188 142 641 3 1 643 DFQD0BWP7T $T=422120 429400 0 0 $X=421830 $Y=429165
X1189 142 653 3 1 637 DFQD0BWP7T $T=436120 390200 1 180 $X=425190 $Y=389965
X1190 142 252 3 1 657 DFQD0BWP7T $T=429400 382360 1 0 $X=429110 $Y=378150
X1191 142 655 3 1 263 DFQD0BWP7T $T=432760 405880 0 0 $X=432470 $Y=405645
X1192 333 3 1 297 304 329 NR3D0BWP7T $T=174040 445080 0 180 $X=170950 $Y=440870
X1193 337 3 1 302 304 29 NR3D0BWP7T $T=174040 476440 1 0 $X=173750 $Y=472230
X1194 570 1 190 192 575 3 AOI21D2BWP7T $T=366680 468600 0 0 $X=366390 $Y=468365
X1195 312 310 306 300 3 1 AOI21D0BWP7T $T=163400 405880 1 180 $X=160310 $Y=405645
X1196 296 331 333 329 3 1 AOI21D0BWP7T $T=172360 437240 1 0 $X=172070 $Y=433030
X1197 25 335 337 29 3 1 AOI21D0BWP7T $T=172920 484280 1 0 $X=172630 $Y=480070
X1198 438 449 443 423 3 1 AOI21D0BWP7T $T=269240 437240 1 180 $X=266150 $Y=437005
X1199 409 3 1 410 BUFFD0BWP7T $T=240680 374520 0 0 $X=240390 $Y=374285
X1200 48 69 3 1 395 AN2D1BWP7T $T=230040 374520 1 180 $X=226950 $Y=374285
X1201 48 101 3 1 419 AN2D1BWP7T $T=259720 429400 1 180 $X=256630 $Y=429165
X1202 111 101 3 1 413 AN2D1BWP7T $T=272040 429400 1 180 $X=268950 $Y=429165
X1203 115 101 3 1 418 AN2D1BWP7T $T=274840 429400 1 180 $X=271750 $Y=429165
X1204 458 102 3 1 113 AN2D1BWP7T $T=276520 366680 0 180 $X=273430 $Y=362470
X1205 96 101 3 1 427 AN2D1BWP7T $T=273720 429400 1 0 $X=273430 $Y=425190
X1206 458 114 3 1 532 AN2D1BWP7T $T=326360 413720 0 0 $X=326070 $Y=413485
X1207 559 454 3 1 562 AN2D1BWP7T $T=350440 452920 1 0 $X=350150 $Y=448710
X1208 559 101 3 1 171 AN2D1BWP7T $T=354360 452920 1 180 $X=351270 $Y=452685
X1209 563 101 3 1 176 AN2D1BWP7T $T=360520 437240 1 180 $X=357430 $Y=437005
X1210 212 101 3 1 584 AN2D1BWP7T $T=395240 429400 1 180 $X=392150 $Y=429165
X1211 231 146 3 1 225 AN2D1BWP7T $T=411480 358840 1 180 $X=408390 $Y=358605
X1212 234 101 3 1 597 AN2D1BWP7T $T=414280 421560 0 180 $X=411190 $Y=417350
X1213 256 101 3 1 596 AN2D1BWP7T $T=433320 437240 1 180 $X=430230 $Y=437005
X1214 261 202 3 1 659 AN2D1BWP7T $T=440600 445080 1 0 $X=440310 $Y=440870
X1215 261 101 3 1 269 AN2D1BWP7T $T=444520 437240 1 180 $X=441430 $Y=437005
X1216 358 375 357 1 3 382 XOR3D0BWP7T $T=209320 405880 1 0 $X=209030 $Y=401670
X1217 463 445 401 1 3 136 XOR3D0BWP7T $T=295000 374520 1 0 $X=294710 $Y=370310
X1218 341 310 313 1 3 350 XNR3D0BWP7T $T=192520 421560 0 180 $X=182710 $Y=417350
X1219 376 407 389 1 3 421 XNR3D0BWP7T $T=249640 413720 0 0 $X=249350 $Y=413485
X1220 436 449 403 1 3 461 XNR3D0BWP7T $T=282680 437240 0 0 $X=282390 $Y=437005
X1221 503 502 515 1 3 519 XNR3D0BWP7T $T=309000 390200 1 0 $X=308710 $Y=385990
X1222 40 42 3 350 1 354 41 OAI22D1BWP7T $T=186360 398040 1 0 $X=186070 $Y=393830
X1223 50 44 3 368 367 1 IOA21D0BWP7T $T=206520 390200 0 180 $X=202870 $Y=385990
X1224 376 389 3 394 416 1 IOA21D0BWP7T $T=248520 429400 0 180 $X=244870 $Y=425190
X1225 95 98 3 104 424 1 IOA21D0BWP7T $T=264200 476440 0 180 $X=260550 $Y=472230
X1226 118 491 3 473 474 1 IOA21D0BWP7T $T=305080 468600 0 180 $X=301430 $Y=464390
X1227 503 515 3 541 528 1 IOA21D0BWP7T $T=328040 398040 0 0 $X=327750 $Y=397805
X1228 469 3 124 117 1 466 474 OAI211D0BWP7T $T=288840 468600 1 0 $X=288550 $Y=464390
X1229 44 71 380 28 3 1 397 AO22D0BWP7T $T=245160 413720 1 180 $X=240390 $Y=413485
X1230 116 124 120 118 3 1 396 AO22D0BWP7T $T=287160 484280 0 180 $X=282390 $Y=480070
X1231 147 124 496 118 3 1 510 AO22D0BWP7T $T=326360 366680 0 0 $X=326070 $Y=366445
X1232 161 124 543 118 3 1 545 AO22D0BWP7T $T=333080 374520 1 0 $X=332790 $Y=370310
X1233 436 403 439 448 3 1 MAOI222D2BWP7T $T=261960 421560 0 0 $X=261670 $Y=421325
X1234 189 194 196 199 3 1 MAOI222D2BWP7T $T=367800 484280 1 0 $X=367510 $Y=480070
X1235 5 293 3 1 9 DFQD1BWP7T $T=156680 390200 1 0 $X=156390 $Y=385990
X1236 5 18 3 1 345 DFQD1BWP7T $T=168440 390200 1 0 $X=168150 $Y=385990
X1237 5 37 3 1 27 DFQD1BWP7T $T=181880 390200 1 0 $X=181590 $Y=385990
X1238 5 49 3 1 38 DFQD1BWP7T $T=209320 382360 1 180 $X=198390 $Y=382125
X1239 5 351 3 1 34 DFQD1BWP7T $T=209320 398040 1 180 $X=198390 $Y=397805
X1240 61 383 3 1 52 DFQD1BWP7T $T=219400 413720 0 180 $X=208470 $Y=409510
X1241 5 354 3 1 64 DFQD1BWP7T $T=211560 390200 0 0 $X=211270 $Y=389965
X1242 5 68 3 1 63 DFQD1BWP7T $T=231720 382360 0 180 $X=220790 $Y=378150
X1243 5 76 3 1 392 DFQD1BWP7T $T=233960 398040 0 180 $X=223030 $Y=393830
X1244 61 397 3 1 83 DFQD1BWP7T $T=223880 460760 1 0 $X=223590 $Y=456550
X1245 61 410 3 1 74 DFQD1BWP7T $T=240680 421560 0 0 $X=240390 $Y=421325
X1246 61 412 3 1 70 DFQD1BWP7T $T=240680 452920 1 0 $X=240390 $Y=448710
X1247 61 414 3 1 91 DFQD1BWP7T $T=241240 460760 0 0 $X=240950 $Y=460525
X1248 61 415 3 1 90 DFQD1BWP7T $T=241240 476440 1 0 $X=240950 $Y=472230
X1249 5 422 3 1 69 DFQD1BWP7T $T=253560 382360 0 180 $X=242630 $Y=378150
X1250 61 430 3 1 94 DFQD1BWP7T $T=263640 468600 0 180 $X=252710 $Y=464390
X1251 5 129 3 1 450 DFQD1BWP7T $T=293320 358840 1 180 $X=282390 $Y=358605
X1252 61 468 3 1 434 DFQD1BWP7T $T=293880 374520 1 180 $X=282950 $Y=374285
X1253 61 467 3 1 132 DFQD1BWP7T $T=303960 468600 1 180 $X=293030 $Y=468365
X1254 142 538 3 1 455 DFQD1BWP7T $T=346520 358840 1 180 $X=335590 $Y=358605
X1255 142 531 3 1 535 DFQD1BWP7T $T=349880 374520 0 180 $X=338950 $Y=370310
X1256 61 169 3 1 178 DFQD1BWP7T $T=348200 468600 1 0 $X=347910 $Y=464390
X1257 142 566 3 1 559 DFQD1BWP7T $T=360520 382360 1 180 $X=349590 $Y=382125
X1258 142 197 3 1 563 DFQD1BWP7T $T=377320 382360 1 180 $X=366390 $Y=382125
X1259 142 581 3 1 191 DFQD1BWP7T $T=379000 358840 1 180 $X=368070 $Y=358605
X1260 142 584 3 1 193 DFQD1BWP7T $T=380680 421560 0 180 $X=369750 $Y=417350
X1261 142 621 3 1 202 DFQD1BWP7T $T=408680 429400 0 0 $X=408390 $Y=429165
X1262 142 658 3 1 223 DFQD1BWP7T $T=443960 421560 1 180 $X=433030 $Y=421325
X1263 44 43 3 1 352 351 41 MOAI22D0BWP7T $T=190840 366680 1 180 $X=186630 $Y=366445
X1264 44 56 3 1 382 383 41 MOAI22D0BWP7T $T=213240 382360 0 0 $X=212950 $Y=382125
X1265 71 406 3 1 40 409 85 MOAI22D0BWP7T $T=246840 374520 1 180 $X=242630 $Y=374285
X1266 118 434 3 1 121 467 119 MOAI22D0BWP7T $T=282680 468600 0 0 $X=282390 $Y=468365
X1267 118 128 3 1 456 468 119 MOAI22D0BWP7T $T=289960 366680 0 180 $X=285750 $Y=362470
X1268 118 450 3 1 133 415 119 MOAI22D0BWP7T $T=297240 476440 1 180 $X=293030 $Y=476205
X1269 118 187 3 1 119 567 560 MOAI22D0BWP7T $T=366680 398040 1 0 $X=366390 $Y=393830
X1270 340 364 51 366 374 3 1 XNR4D0BWP7T $T=198680 374520 1 0 $X=198390 $Y=370310
X1271 53 314 388 390 66 3 1 XNR4D0BWP7T $T=209880 476440 1 0 $X=209590 $Y=472230
X1272 542 550 555 551 523 3 1 XNR4D0BWP7T $T=334760 452920 1 0 $X=334470 $Y=448710
X1273 555 564 560 549 536 3 1 XNR4D0BWP7T $T=359400 413720 0 180 $X=346230 $Y=409510
X1274 275 267 259 258 648 3 1 XNR4D0BWP7T $T=444520 452920 1 180 $X=431350 $Y=452685
X1275 40 3 89 412 41 421 1 OAI22D2BWP7T $T=244040 398040 0 0 $X=243750 $Y=397805
X1276 373 339 366 343 47 3 1 XOR4D0BWP7T $T=211560 358840 1 180 $X=198390 $Y=358605
X1277 78 399 390 378 379 3 1 XOR4D0BWP7T $T=232840 445080 1 180 $X=219670 $Y=444845
X1278 93 420 88 86 408 3 1 XOR4D0BWP7T $T=253560 366680 0 180 $X=240390 $Y=362470
X1279 544 488 536 533 145 3 1 XOR4D0BWP7T $T=337560 429400 0 180 $X=324390 $Y=425190
X1280 526 534 551 524 554 3 1 XOR4D0BWP7T $T=330840 437240 0 0 $X=330550 $Y=437005
X1281 556 553 549 547 521 3 1 XOR4D0BWP7T $T=346520 413720 0 180 $X=333350 $Y=409510
X1282 7 3 1 295 CKND1BWP7T $T=158920 468600 0 0 $X=158630 $Y=468365
X1283 345 12 3 1 BUFFD1P5BWP7T $T=179080 390200 1 0 $X=178790 $Y=385990
X1284 392 31 3 1 BUFFD1P5BWP7T $T=220520 398040 1 0 $X=220230 $Y=393830
X1285 262 188 1 3 CKND2BWP7T $T=438920 429400 1 180 $X=436390 $Y=429165
X1286 294 3 1 7 CKBD1BWP7T $T=158360 445080 0 0 $X=158070 $Y=444845
X1287 298 3 1 292 CKBD1BWP7T $T=159480 398040 0 0 $X=159190 $Y=397805
X1288 330 3 1 22 CKBD1BWP7T $T=171240 405880 1 0 $X=170950 $Y=401670
X1289 321 3 1 23 CKBD1BWP7T $T=172920 413720 0 0 $X=172630 $Y=413485
X1290 417 3 1 87 CKBD1BWP7T $T=246840 484280 0 180 $X=244310 $Y=480070
X1291 440 3 1 107 CKBD1BWP7T $T=267000 476440 1 0 $X=266710 $Y=472230
X1292 149 3 1 471 CKBD1BWP7T $T=328600 382360 1 180 $X=326070 $Y=382125
X1293 164 3 1 470 CKBD1BWP7T $T=339240 468600 1 0 $X=338950 $Y=464390
X1294 170 3 1 454 CKBD1BWP7T $T=352120 460760 1 180 $X=349590 $Y=460525
X1295 558 3 1 529 CKBD1BWP7T $T=354360 398040 1 180 $X=351830 $Y=397805
X1296 573 3 1 458 CKBD1BWP7T $T=370600 421560 1 180 $X=368070 $Y=421325
X1297 557 3 1 145 CKBD1BWP7T $T=370600 429400 1 180 $X=368070 $Y=429165
X1298 552 3 1 153 CKBD1BWP7T $T=382920 429400 0 180 $X=380390 $Y=425190
X1299 583 3 1 156 CKBD1BWP7T $T=392440 382360 0 180 $X=389910 $Y=378150
X1300 588 647 648 243 650 3 1 OAI31D1BWP7T $T=426040 452920 1 0 $X=425750 $Y=448710
X1301 55 28 340 1 3 384 OA21D0BWP7T $T=213240 358840 0 0 $X=212950 $Y=358605
X1302 153 539 542 1 3 513 OA21D0BWP7T $T=328600 452920 1 0 $X=328310 $Y=448710
X1303 251 644 249 1 3 248 OA21D0BWP7T $T=429400 476440 1 180 $X=425750 $Y=476205
X1304 227 616 219 614 611 1 3 AOI22D0BWP7T $T=402520 398040 1 180 $X=398870 $Y=397805
X1305 233 612 219 594 618 1 3 AOI22D0BWP7T $T=412040 374520 1 180 $X=408390 $Y=374285
X1306 227 622 219 608 594 1 3 AOI22D0BWP7T $T=414840 390200 1 180 $X=411190 $Y=389965
X1307 230 624 219 615 237 1 3 AOI22D0BWP7T $T=413720 366680 0 0 $X=413430 $Y=366445
X1308 608 628 629 219 228 1 3 AOI22D0BWP7T $T=413720 405880 1 0 $X=413430 $Y=401670
X1309 233 627 219 611 615 1 3 AOI22D0BWP7T $T=417640 382360 1 180 $X=413990 $Y=382125
X1310 230 236 219 618 238 1 3 AOI22D0BWP7T $T=415960 358840 0 0 $X=415670 $Y=358605
X1311 614 623 202 219 228 1 3 AOI22D0BWP7T $T=417080 413720 1 0 $X=416790 $Y=409510
X1312 227 638 219 634 637 1 3 AOI22D0BWP7T $T=419880 390200 0 0 $X=419590 $Y=389965
X1313 233 639 219 637 630 1 3 AOI22D0BWP7T $T=424360 382360 1 180 $X=420710 $Y=382125
X1314 230 642 219 630 633 1 3 AOI22D0BWP7T $T=426040 374520 0 180 $X=422390 $Y=370310
X1315 250 651 219 633 253 1 3 AOI22D0BWP7T $T=428840 366680 1 0 $X=428550 $Y=362470
X1316 634 645 643 219 228 1 3 AOI22D0BWP7T $T=434440 413720 0 0 $X=434150 $Y=413485
X1317 227 656 219 263 266 1 3 AOI22D0BWP7T $T=437800 398040 0 0 $X=437510 $Y=397805
X1318 233 264 219 266 657 1 3 AOI22D0BWP7T $T=439480 390200 1 0 $X=439190 $Y=385990
X1319 230 265 219 657 272 1 3 AOI22D0BWP7T $T=440040 374520 1 0 $X=439750 $Y=370310
X1320 268 270 219 253 276 1 3 AOI22D0BWP7T $T=441160 366680 1 0 $X=440870 $Y=362470
X1321 3 1 ICV_76 $T=155000 358840 0 0 $X=154710 $Y=358605
X1322 3 1 ICV_76 $T=155000 366680 0 0 $X=154710 $Y=366445
X1323 3 1 ICV_76 $T=155000 476440 0 0 $X=154710 $Y=476205
X1324 3 1 ICV_76 $T=197000 366680 1 0 $X=196710 $Y=362470
X1325 3 1 ICV_76 $T=197000 374520 0 0 $X=196710 $Y=374285
X1326 3 1 ICV_76 $T=197000 398040 1 0 $X=196710 $Y=393830
X1327 3 1 ICV_76 $T=197000 429400 1 0 $X=196710 $Y=425190
X1328 3 1 ICV_76 $T=197000 429400 0 0 $X=196710 $Y=429165
X1329 3 1 ICV_76 $T=239000 405880 1 0 $X=238710 $Y=401670
X1330 3 1 ICV_76 $T=239000 413720 1 0 $X=238710 $Y=409510
X1331 3 1 ICV_76 $T=239000 445080 0 0 $X=238710 $Y=444845
X1332 3 1 ICV_76 $T=281000 413720 1 0 $X=280710 $Y=409510
X1333 3 1 ICV_76 $T=365000 390200 1 0 $X=364710 $Y=385990
X1334 3 1 ICV_76 $T=365000 398040 0 0 $X=364710 $Y=397805
X1335 3 1 ICV_76 $T=365000 460760 1 0 $X=364710 $Y=456550
X1336 3 1 ICV_76 $T=407000 382360 1 0 $X=406710 $Y=378150
X1337 3 1 ICV_76 $T=407000 390200 1 0 $X=406710 $Y=385990
X1338 3 1 ICV_76 $T=407000 413720 0 0 $X=406710 $Y=413485
X1339 3 1 ICV_76 $T=407000 429400 1 0 $X=406710 $Y=425190
X1340 3 1 ICV_41 $T=156120 421560 0 0 $X=155830 $Y=421325
X1341 3 1 ICV_41 $T=198120 390200 0 0 $X=197830 $Y=389965
X1342 3 1 ICV_41 $T=224440 390200 1 0 $X=224150 $Y=385990
X1343 3 1 ICV_41 $T=240120 374520 1 0 $X=239830 $Y=370310
X1344 3 1 ICV_41 $T=240120 437240 0 0 $X=239830 $Y=437005
X1345 3 1 ICV_41 $T=307880 421560 1 0 $X=307590 $Y=417350
X1346 3 1 ICV_41 $T=307880 452920 0 0 $X=307590 $Y=452685
X1347 3 1 ICV_41 $T=307880 468600 1 0 $X=307590 $Y=464390
X1348 3 1 ICV_41 $T=309560 476440 0 0 $X=309270 $Y=476205
X1349 3 1 ICV_41 $T=324120 366680 1 0 $X=323830 $Y=362470
X1350 3 1 ICV_41 $T=344280 437240 1 0 $X=343990 $Y=433030
X1351 3 1 ICV_41 $T=349880 374520 1 0 $X=349590 $Y=370310
X1352 3 1 ICV_41 $T=350440 429400 1 0 $X=350150 $Y=425190
X1353 3 1 ICV_41 $T=366120 429400 1 0 $X=365830 $Y=425190
X1354 3 1 ICV_41 $T=375080 484280 1 0 $X=374790 $Y=480070
X1355 3 1 ICV_41 $T=377320 374520 1 0 $X=377030 $Y=370310
X1356 3 1 ICV_41 $T=392440 382360 1 0 $X=392150 $Y=378150
X1357 3 1 ICV_41 $T=392440 421560 0 0 $X=392150 $Y=421325
X1358 3 1 ICV_41 $T=408120 374520 1 0 $X=407830 $Y=370310
X1359 3 1 ICV_37 $T=156120 398040 0 0 $X=155830 $Y=397805
X1360 3 1 ICV_37 $T=156120 413720 0 0 $X=155830 $Y=413485
X1361 3 1 ICV_37 $T=156120 476440 1 0 $X=155830 $Y=472230
X1362 3 1 ICV_37 $T=163400 405880 0 0 $X=163110 $Y=405645
X1363 3 1 ICV_37 $T=165080 445080 0 0 $X=164790 $Y=444845
X1364 3 1 ICV_37 $T=167320 421560 1 0 $X=167030 $Y=417350
X1365 3 1 ICV_37 $T=172360 421560 1 0 $X=172070 $Y=417350
X1366 3 1 ICV_37 $T=193640 429400 1 0 $X=193350 $Y=425190
X1367 3 1 ICV_37 $T=193640 484280 1 0 $X=193350 $Y=480070
X1368 3 1 ICV_37 $T=207080 366680 0 0 $X=206790 $Y=366445
X1369 3 1 ICV_37 $T=209320 382360 0 0 $X=209030 $Y=382125
X1370 3 1 ICV_37 $T=224440 460760 0 0 $X=224150 $Y=460525
X1371 3 1 ICV_37 $T=235640 429400 0 0 $X=235350 $Y=429165
X1372 3 1 ICV_37 $T=249080 390200 1 0 $X=248790 $Y=385990
X1373 3 1 ICV_37 $T=260280 390200 0 0 $X=259990 $Y=389965
X1374 3 1 ICV_37 $T=282120 374520 1 0 $X=281830 $Y=370310
X1375 3 1 ICV_37 $T=282120 452920 1 0 $X=281830 $Y=448710
X1376 3 1 ICV_37 $T=291080 429400 0 0 $X=290790 $Y=429165
X1377 3 1 ICV_37 $T=324120 358840 0 0 $X=323830 $Y=358605
X1378 3 1 ICV_37 $T=324120 398040 1 0 $X=323830 $Y=393830
X1379 3 1 ICV_37 $T=324120 460760 1 0 $X=323830 $Y=456550
X1380 3 1 ICV_37 $T=343720 437240 0 0 $X=343430 $Y=437005
X1381 3 1 ICV_37 $T=375080 366680 0 0 $X=374790 $Y=366445
X1382 3 1 ICV_37 $T=377320 445080 1 0 $X=377030 $Y=440870
X1383 3 1 ICV_37 $T=392440 413720 1 0 $X=392150 $Y=409510
X1384 3 1 ICV_37 $T=403640 445080 1 0 $X=403350 $Y=440870
X1385 3 1 ICV_37 $T=408120 421560 1 0 $X=407830 $Y=417350
X1386 3 1 ICV_37 $T=408120 445080 0 0 $X=407830 $Y=444845
X1387 3 1 ICV_37 $T=412600 398040 0 0 $X=412310 $Y=397805
X1388 3 1 ICV_37 $T=417640 382360 0 0 $X=417350 $Y=382125
X1389 3 1 ICV_37 $T=426040 382360 1 0 $X=425750 $Y=378150
X1390 3 1 ICV_37 $T=427160 437240 0 0 $X=426870 $Y=437005
X1391 3 1 ICV_37 $T=428840 445080 1 0 $X=428550 $Y=440870
X1392 3 1 ICV_37 $T=436120 390200 1 0 $X=435830 $Y=385990
X1393 3 1 ICV_37 $T=437800 413720 0 0 $X=437510 $Y=413485
X1394 3 1 ICV_37 $T=445640 484280 1 0 $X=445350 $Y=480070
X1395 3 1 ICV_43 $T=156120 468600 0 0 $X=155830 $Y=468365
X1396 3 1 ICV_43 $T=170680 398040 0 0 $X=170390 $Y=397805
X1397 3 1 ICV_43 $T=207080 476440 1 0 $X=206790 $Y=472230
X1398 3 1 ICV_43 $T=217720 421560 1 0 $X=217430 $Y=417350
X1399 3 1 ICV_43 $T=225000 429400 0 0 $X=224710 $Y=429165
X1400 3 1 ICV_43 $T=225000 476440 0 0 $X=224710 $Y=476205
X1401 3 1 ICV_43 $T=240120 382360 1 0 $X=239830 $Y=378150
X1402 3 1 ICV_43 $T=264200 476440 1 0 $X=263910 $Y=472230
X1403 3 1 ICV_43 $T=266440 405880 1 0 $X=266150 $Y=401670
X1404 3 1 ICV_43 $T=269240 405880 0 0 $X=268950 $Y=405645
X1405 3 1 ICV_43 $T=282120 468600 1 0 $X=281830 $Y=464390
X1406 3 1 ICV_43 $T=291080 398040 0 0 $X=290790 $Y=397805
X1407 3 1 ICV_43 $T=307880 366680 1 0 $X=307590 $Y=362470
X1408 3 1 ICV_43 $T=331400 398040 0 0 $X=331110 $Y=397805
X1409 3 1 ICV_43 $T=331960 452920 1 0 $X=331670 $Y=448710
X1410 3 1 ICV_43 $T=347640 452920 1 0 $X=347350 $Y=448710
X1411 3 1 ICV_43 $T=355480 358840 0 0 $X=355190 $Y=358605
X1412 3 1 ICV_43 $T=385160 445080 1 0 $X=384870 $Y=440870
X1413 3 1 ICV_43 $T=391880 429400 1 0 $X=391590 $Y=425190
X1414 3 1 ICV_43 $T=394680 445080 1 0 $X=394390 $Y=440870
X1415 3 1 ICV_43 $T=420440 413720 1 0 $X=420150 $Y=409510
X1416 3 1 ICV_43 $T=426040 366680 1 0 $X=425750 $Y=362470
X1417 3 1 ICV_43 $T=446200 445080 0 0 $X=445910 $Y=444845
X1418 3 1 ICV_52 $T=193080 413720 0 0 $X=192790 $Y=413485
X1419 3 1 ICV_52 $T=235080 382360 0 0 $X=234790 $Y=382125
X1420 3 1 ICV_52 $T=240120 398040 0 0 $X=239830 $Y=397805
X1421 3 1 ICV_52 $T=249080 358840 0 0 $X=248790 $Y=358605
X1422 3 1 ICV_52 $T=249080 452920 0 0 $X=248790 $Y=452685
X1423 3 1 ICV_52 $T=249080 468600 1 0 $X=248790 $Y=464390
X1424 3 1 ICV_52 $T=255800 452920 1 0 $X=255510 $Y=448710
X1425 3 1 ICV_52 $T=257480 437240 0 0 $X=257190 $Y=437005
X1426 3 1 ICV_52 $T=258040 413720 1 0 $X=257750 $Y=409510
X1427 3 1 ICV_52 $T=291080 398040 1 0 $X=290790 $Y=393830
X1428 3 1 ICV_52 $T=303960 468600 0 0 $X=303670 $Y=468365
X1429 3 1 ICV_52 $T=319080 437240 0 0 $X=318790 $Y=437005
X1430 3 1 ICV_52 $T=324120 468600 1 0 $X=323830 $Y=464390
X1431 3 1 ICV_52 $T=361080 390200 1 0 $X=360790 $Y=385990
X1432 3 1 ICV_52 $T=366120 421560 1 0 $X=365830 $Y=417350
X1433 3 1 ICV_52 $T=384040 398040 0 0 $X=383750 $Y=397805
X1434 3 1 ICV_52 $T=387960 358840 0 0 $X=387670 $Y=358605
X1435 3 1 ICV_52 $T=395240 452920 0 0 $X=394950 $Y=452685
X1436 3 1 ICV_52 $T=417080 405880 1 0 $X=416790 $Y=401670
X1437 3 1 ICV_52 $T=417080 460760 0 0 $X=416790 $Y=460525
X1438 3 1 ICV_52 $T=427720 452920 0 0 $X=427430 $Y=452685
X1439 3 1 ICV_52 $T=427720 468600 0 0 $X=427430 $Y=468365
X1440 3 1 ICV_52 $T=436120 374520 1 0 $X=435830 $Y=370310
X1441 3 1 ICV_52 $T=445080 374520 0 0 $X=444790 $Y=374285
X1442 3 1 ICV_52 $T=445080 390200 0 0 $X=444790 $Y=389965
X1443 3 1 ICV_54 $T=169000 429400 0 0 $X=168710 $Y=429165
X1444 3 1 ICV_54 $T=174040 476440 0 0 $X=173750 $Y=476205
X1445 3 1 ICV_54 $T=191400 405880 1 0 $X=191110 $Y=401670
X1446 3 1 ICV_54 $T=191400 405880 0 0 $X=191110 $Y=405645
X1447 3 1 ICV_54 $T=216040 366680 1 0 $X=215750 $Y=362470
X1448 3 1 ICV_54 $T=275400 405880 0 0 $X=275110 $Y=405645
X1449 3 1 ICV_54 $T=275400 413720 1 0 $X=275110 $Y=409510
X1450 3 1 ICV_54 $T=275400 452920 1 0 $X=275110 $Y=448710
X1451 3 1 ICV_54 $T=293320 358840 0 0 $X=293030 $Y=358605
X1452 3 1 ICV_54 $T=300040 460760 1 0 $X=299750 $Y=456550
X1453 3 1 ICV_54 $T=330280 358840 0 0 $X=329990 $Y=358605
X1454 3 1 ICV_54 $T=359400 413720 1 0 $X=359110 $Y=409510
X1455 3 1 ICV_54 $T=384040 390200 1 0 $X=383750 $Y=385990
X1456 3 1 ICV_54 $T=401400 452920 0 0 $X=401110 $Y=452685
X1457 3 1 ICV_54 $T=401400 468600 1 0 $X=401110 $Y=464390
X1458 3 1 ICV_54 $T=408120 405880 1 0 $X=407830 $Y=401670
X1459 3 1 ICV_54 $T=443400 374520 1 0 $X=443110 $Y=370310
X1460 3 1 ICV_54 $T=443400 405880 0 0 $X=443110 $Y=405645
X1461 174 1 188 185 3 NR2XD0BWP7T $T=368920 452920 0 180 $X=366390 $Y=448710
X1462 119 124 3 1 INVD2P5BWP7T $T=298920 358840 0 0 $X=298630 $Y=358605
X1463 143 3 1 100 BUFFD3BWP7T $T=317400 484280 0 180 $X=313190 $Y=480070
X1464 450 446 3 1 451 453 IAO21D0BWP7T $T=269240 405880 1 0 $X=268950 $Y=401670
X1465 116 400 3 1 464 465 IAO21D0BWP7T $T=282680 413720 0 0 $X=282390 $Y=413485
X1466 492 509 3 1 505 499 IAO21D0BWP7T $T=311240 468600 0 0 $X=310950 $Y=468365
X1467 178 599 3 1 598 585 IAO21D0BWP7T $T=392440 468600 0 180 $X=388790 $Y=464390
X1468 215 613 3 1 222 604 IAO21D0BWP7T $T=399160 468600 0 0 $X=398870 $Y=468365
X1469 112 455 450 1 3 451 AN3D1BWP7T $T=275400 405880 1 180 $X=271750 $Y=405645
X1470 112 471 116 1 3 464 AN3D1BWP7T $T=289960 421560 0 180 $X=286310 $Y=417350
X1471 112 529 492 1 3 505 AN3D1BWP7T $T=329160 468600 1 180 $X=325510 $Y=468365
X1472 207 211 178 1 3 598 AN3D1BWP7T $T=395800 468600 0 180 $X=392150 $Y=464390
X1473 207 223 215 1 3 222 AN3D1BWP7T $T=424360 484280 0 180 $X=420710 $Y=480070
X1474 207 629 246 1 3 244 AN3D1BWP7T $T=427720 484280 0 180 $X=424070 $Y=480070
X1475 61 368 75 3 1 DFQD2BWP7T $T=220520 421560 1 0 $X=220230 $Y=417350
X1477 3 1 ICV_80 $T=407000 468600 1 0 $X=406710 $Y=464390
X1478 3 1 ICV_64 $T=191960 445080 1 0 $X=191670 $Y=440870
X1479 3 1 ICV_64 $T=191960 445080 0 0 $X=191670 $Y=444845
X1480 3 1 ICV_64 $T=191960 452920 1 0 $X=191670 $Y=448710
X1481 3 1 ICV_64 $T=233960 398040 1 0 $X=233670 $Y=393830
X1482 3 1 ICV_64 $T=233960 437240 0 0 $X=233670 $Y=437005
X1483 3 1 ICV_64 $T=233960 445080 1 0 $X=233670 $Y=440870
X1484 3 1 ICV_64 $T=233960 468600 1 0 $X=233670 $Y=464390
X1485 3 1 ICV_64 $T=233960 468600 0 0 $X=233670 $Y=468365
X1486 3 1 ICV_64 $T=275960 382360 0 0 $X=275670 $Y=382125
X1487 3 1 ICV_64 $T=275960 398040 1 0 $X=275670 $Y=393830
X1488 3 1 ICV_64 $T=275960 445080 1 0 $X=275670 $Y=440870
X1489 3 1 ICV_64 $T=275960 468600 1 0 $X=275670 $Y=464390
X1490 3 1 ICV_64 $T=275960 468600 0 0 $X=275670 $Y=468365
X1491 3 1 ICV_64 $T=317960 366680 0 0 $X=317670 $Y=366445
X1492 3 1 ICV_64 $T=317960 374520 0 0 $X=317670 $Y=374285
X1493 3 1 ICV_64 $T=317960 382360 0 0 $X=317670 $Y=382125
X1494 3 1 ICV_64 $T=317960 421560 0 0 $X=317670 $Y=421325
X1495 3 1 ICV_64 $T=317960 437240 1 0 $X=317670 $Y=433030
X1496 3 1 ICV_64 $T=317960 476440 1 0 $X=317670 $Y=472230
X1497 3 1 ICV_64 $T=359960 405880 0 0 $X=359670 $Y=405645
X1498 3 1 ICV_64 $T=359960 476440 1 0 $X=359670 $Y=472230
X1499 3 1 ICV_64 $T=401960 374520 0 0 $X=401670 $Y=374285
X1500 3 1 ICV_64 $T=401960 405880 1 0 $X=401670 $Y=401670
X1501 3 1 ICV_64 $T=401960 445080 0 0 $X=401670 $Y=444845
X1502 3 1 ICV_64 $T=401960 460760 1 0 $X=401670 $Y=456550
X1503 3 1 ICV_64 $T=401960 476440 1 0 $X=401670 $Y=472230
X1504 3 1 ICV_81 $T=155000 374520 1 0 $X=154710 $Y=370310
X1505 3 1 ICV_81 $T=155000 382360 1 0 $X=154710 $Y=378150
X1506 3 1 ICV_81 $T=155000 390200 0 0 $X=154710 $Y=389965
X1507 3 1 ICV_81 $T=155000 413720 1 0 $X=154710 $Y=409510
X1508 3 1 ICV_81 $T=155000 468600 1 0 $X=154710 $Y=464390
X1509 3 1 ICV_81 $T=197000 413720 0 0 $X=196710 $Y=413485
X1510 3 1 ICV_81 $T=197000 452920 0 0 $X=196710 $Y=452685
X1511 3 1 ICV_81 $T=197000 484280 1 0 $X=196710 $Y=480070
X1512 3 1 ICV_81 $T=239000 366680 0 0 $X=238710 $Y=366445
X1513 3 1 ICV_81 $T=239000 460760 1 0 $X=238710 $Y=456550
X1514 3 1 ICV_81 $T=239000 476440 0 0 $X=238710 $Y=476205
X1515 3 1 ICV_81 $T=281000 405880 0 0 $X=280710 $Y=405645
X1516 3 1 ICV_81 $T=281000 460760 0 0 $X=280710 $Y=460525
X1517 3 1 ICV_81 $T=323000 405880 1 0 $X=322710 $Y=401670
X1518 3 1 ICV_81 $T=323000 421560 1 0 $X=322710 $Y=417350
X1519 3 1 ICV_81 $T=323000 429400 0 0 $X=322710 $Y=429165
X1520 3 1 ICV_81 $T=365000 366680 1 0 $X=364710 $Y=362470
X1521 3 1 ICV_81 $T=365000 390200 0 0 $X=364710 $Y=389965
X1522 3 1 ICV_69 $T=155000 429400 1 0 $X=154710 $Y=425190
X1523 3 1 ICV_69 $T=155000 437240 0 0 $X=154710 $Y=437005
X1524 3 1 ICV_69 $T=197000 366680 0 0 $X=196710 $Y=366445
X1525 3 1 ICV_69 $T=197000 405880 1 0 $X=196710 $Y=401670
X1526 3 1 ICV_69 $T=197000 421560 0 0 $X=196710 $Y=421325
X1527 3 1 ICV_69 $T=197000 476440 1 0 $X=196710 $Y=472230
X1528 3 1 ICV_69 $T=239000 358840 0 0 $X=238710 $Y=358605
X1529 3 1 ICV_69 $T=239000 390200 1 0 $X=238710 $Y=385990
X1530 3 1 ICV_69 $T=239000 429400 0 0 $X=238710 $Y=429165
X1531 3 1 ICV_69 $T=281000 390200 1 0 $X=280710 $Y=385990
X1532 3 1 ICV_69 $T=281000 398040 0 0 $X=280710 $Y=397805
X1533 3 1 ICV_69 $T=281000 429400 0 0 $X=280710 $Y=429165
X1534 3 1 ICV_69 $T=365000 366680 0 0 $X=364710 $Y=366445
X1535 3 1 ICV_69 $T=365000 452920 0 0 $X=364710 $Y=452685
X1536 3 1 ICV_69 $T=407000 437240 0 0 $X=406710 $Y=437005
X1537 3 1 ICV_69 $T=407000 452920 1 0 $X=406710 $Y=448710
X1538 3 1 ICV_69 $T=407000 452920 0 0 $X=406710 $Y=452685
X1539 3 1 ICV_69 $T=407000 460760 0 0 $X=406710 $Y=460525
X1540 3 1 ICV_69 $T=407000 484280 1 0 $X=406710 $Y=480070
X1541 387 3 71 338 1 367 75 OAI211D1BWP7T $T=227800 429400 0 0 $X=227510 $Y=429165
X1542 100 3 102 41 1 ND2D4BWP7T $T=253560 374520 1 0 $X=253270 $Y=370310
X1543 97 1 100 3 44 NR2XD3BWP7T $T=254680 398040 0 0 $X=254390 $Y=397805
X1544 408 44 3 41 414 388 1 MOAI22D1BWP7T $T=266440 413720 0 180 $X=261670 $Y=409510
X1545 118 125 3 119 447 461 1 MOAI22D1BWP7T $T=287720 429400 0 180 $X=282950 $Y=425190
X1546 118 492 3 119 135 134 1 MOAI22D1BWP7T $T=304520 484280 0 180 $X=299750 $Y=480070
X1547 118 160 3 119 537 519 1 MOAI22D1BWP7T $T=333640 390200 0 180 $X=328870 $Y=385990
X1548 119 1 140 525 3 511 508 AOI211D1BWP7T $T=328040 374520 1 180 $X=324390 $Y=374285
X1549 546 1 119 162 3 165 163 AOI211D1BWP7T $T=339240 366680 1 0 $X=338950 $Y=362470
X1550 10 148 514 1 3 NR2D1P5BWP7T $T=328600 437240 1 180 $X=324390 $Y=437005
X1551 172 10 3 1 BUFFD8BWP7T $T=356040 437240 1 180 $X=346790 $Y=437005
.ENDS
***************************************
.SUBCKT IAO21D1BWP7T A1 A2 VDD B ZN VSS
** N=9 EP=6 IP=0 FDC=8
*.SEEDPROM
M0 7 A1 VSS VSS N L=1.8e-07 W=5.7e-07 $X=730 $Y=345 $D=0
M1 VSS A2 7 VSS N L=1.8e-07 W=5.7e-07 $X=1450 $Y=345 $D=0
M2 ZN 7 VSS VSS N L=1.8e-07 W=1e-06 $X=2230 $Y=345 $D=0
M3 VSS B ZN VSS N L=1.8e-07 W=1e-06 $X=2950 $Y=345 $D=0
M4 8 A1 7 VDD P L=1.8e-07 W=8.1e-07 $X=730 $Y=2765 $D=16
M5 VDD A2 8 VDD P L=1.8e-07 W=8.1e-07 $X=1330 $Y=2765 $D=16
M6 9 7 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2230 $Y=2205 $D=16
M7 ZN B 9 VDD P L=1.8e-07 W=1.37e-06 $X=2830 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IOA22D2BWP7T A1 A2 ZN B2 VDD B1 VSS
** N=12 EP=7 IP=0 FDC=14
*.SEEDPROM
M0 9 10 VSS VSS N L=1.8e-07 W=1e-06 $X=660 $Y=345 $D=0
M1 11 A1 9 VSS N L=1.8e-07 W=1e-06 $X=1595 $Y=345 $D=0
M2 VSS A2 11 VSS N L=1.8e-07 W=1e-06 $X=2140 $Y=345 $D=0
M3 ZN 9 VSS VSS N L=1.8e-07 W=1e-06 $X=3235 $Y=345 $D=0
M4 VSS 9 ZN VSS N L=1.8e-07 W=1e-06 $X=3955 $Y=345 $D=0
M5 10 B2 VSS VSS N L=1.8e-07 W=5e-07 $X=4640 $Y=845 $D=0
M6 VSS B1 10 VSS N L=1.8e-07 W=5e-07 $X=5360 $Y=845 $D=0
M7 8 10 9 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M8 VDD A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M9 8 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2070 $Y=2205 $D=16
M10 ZN 9 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3345 $Y=2205 $D=16
M11 VDD 9 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4065 $Y=2205 $D=16
M12 12 B2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4805 $Y=2205 $D=16
M13 10 B1 12 VDD P L=1.8e-07 W=1.37e-06 $X=5360 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INVD10BWP7T I ZN VSS VDD
** N=4 EP=4 IP=0 FDC=20
*.SEEDPROM
M0 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=650 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=1370 $Y=345 $D=0
M2 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=2150 $Y=345 $D=0
M3 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=2870 $Y=345 $D=0
M4 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=3650 $Y=345 $D=0
M5 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=4370 $Y=345 $D=0
M6 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=5150 $Y=345 $D=0
M7 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=5870 $Y=345 $D=0
M8 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=6630 $Y=345 $D=0
M9 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=7350 $Y=345 $D=0
M10 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=650 $Y=2205 $D=16
M11 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1370 $Y=2205 $D=16
M12 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=2150 $Y=2205 $D=16
M13 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=2870 $Y=2205 $D=16
M14 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=3650 $Y=2205 $D=16
M15 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=4370 $Y=2205 $D=16
M16 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=5150 $Y=2205 $D=16
M17 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=5870 $Y=2205 $D=16
M18 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=6630 $Y=2205 $D=16
M19 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=7350 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INR2XD4BWP7T B1 ZN A1 VSS VDD
** N=7 EP=5 IP=0 FDC=32
*.SEEDPROM
M0 ZN B1 VSS VSS N L=1.8e-07 W=5.7e-07 $X=620 $Y=345 $D=0
M1 VSS B1 ZN VSS N L=1.8e-07 W=5.7e-07 $X=1340 $Y=345 $D=0
M2 ZN B1 VSS VSS N L=1.8e-07 W=5.7e-07 $X=2060 $Y=345 $D=0
M3 VSS B1 ZN VSS N L=1.8e-07 W=5.7e-07 $X=2780 $Y=345 $D=0
M4 ZN B1 VSS VSS N L=1.8e-07 W=5.7e-07 $X=3500 $Y=345 $D=0
M5 VSS B1 ZN VSS N L=1.8e-07 W=5.7e-07 $X=4220 $Y=345 $D=0
M6 ZN B1 VSS VSS N L=1.8e-07 W=5.7e-07 $X=4940 $Y=345 $D=0
M7 VSS 7 ZN VSS N L=1.8e-07 W=5.7e-07 $X=5660 $Y=345 $D=0
M8 ZN 7 VSS VSS N L=1.8e-07 W=5.7e-07 $X=6380 $Y=345 $D=0
M9 VSS 7 ZN VSS N L=1.8e-07 W=5.7e-07 $X=7100 $Y=345 $D=0
M10 ZN 7 VSS VSS N L=1.8e-07 W=5.7e-07 $X=7820 $Y=345 $D=0
M11 VSS 7 ZN VSS N L=1.8e-07 W=5.7e-07 $X=8540 $Y=345 $D=0
M12 ZN 7 VSS VSS N L=1.8e-07 W=5.7e-07 $X=9260 $Y=345 $D=0
M13 VSS 7 ZN VSS N L=1.8e-07 W=5.7e-07 $X=9980 $Y=345 $D=0
M14 7 A1 VSS VSS N L=1.8e-07 W=1e-06 $X=11360 $Y=345 $D=0
M15 VSS A1 7 VSS N L=1.8e-07 W=1e-06 $X=12080 $Y=345 $D=0
M16 6 B1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M17 VDD B1 6 VDD P L=1.8e-07 W=1.555e-06 $X=1340 $Y=2020 $D=16
M18 6 B1 VDD VDD P L=1.8e-07 W=1.555e-06 $X=2060 $Y=2020 $D=16
M19 VDD B1 6 VDD P L=1.8e-07 W=1.555e-06 $X=2780 $Y=2020 $D=16
M20 6 B1 VDD VDD P L=1.8e-07 W=1.555e-06 $X=3500 $Y=2020 $D=16
M21 VDD B1 6 VDD P L=1.8e-07 W=1.555e-06 $X=4220 $Y=2020 $D=16
M22 6 B1 VDD VDD P L=1.8e-07 W=1.555e-06 $X=4940 $Y=2020 $D=16
M23 ZN 7 6 VDD P L=1.8e-07 W=1.555e-06 $X=5660 $Y=2020 $D=16
M24 6 7 ZN VDD P L=1.8e-07 W=1.555e-06 $X=6380 $Y=2020 $D=16
M25 ZN 7 6 VDD P L=1.8e-07 W=1.555e-06 $X=7100 $Y=2020 $D=16
M26 6 7 ZN VDD P L=1.8e-07 W=1.555e-06 $X=7820 $Y=2020 $D=16
M27 ZN 7 6 VDD P L=1.8e-07 W=1.555e-06 $X=8540 $Y=2020 $D=16
M28 6 7 ZN VDD P L=1.8e-07 W=1.555e-06 $X=9260 $Y=2020 $D=16
M29 ZN 7 6 VDD P L=1.8e-07 W=1.37e-06 $X=9980 $Y=2205 $D=16
M30 7 A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=11360 $Y=2205 $D=16
M31 VDD A1 7 VDD P L=1.8e-07 W=1.37e-06 $X=12080 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ND3D1BWP7T A3 VSS A2 A1 VDD ZN
** N=8 EP=6 IP=0 FDC=6
*.SEEDPROM
M0 7 A3 VSS VSS N L=1.8e-07 W=1e-06 $X=750 $Y=345 $D=0
M1 8 A2 7 VSS N L=1.8e-07 W=1e-06 $X=1350 $Y=345 $D=0
M2 ZN A1 8 VSS N L=1.8e-07 W=1e-06 $X=1950 $Y=345 $D=0
M3 ZN A3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=750 $Y=2205 $D=16
M4 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1470 $Y=2205 $D=16
M5 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2190 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_79 1 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23
+ 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43
+ 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63
+ 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143
+ 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183
+ 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203
+ 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223
+ 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243
+ 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 262 263
+ 264 265 266 267 268 269
** N=605 EP=266 IP=3984 FDC=10910
*.SEEDPROM
M0 600 129 5 5 N L=1.8e-07 W=1e-06 $X=297540 $Y=594385 $D=0
M1 123 127 600 5 N L=1.8e-07 W=1e-06 $X=298080 $Y=594385 $D=0
M2 601 127 123 5 N L=1.8e-07 W=1e-06 $X=298840 $Y=594385 $D=0
M3 5 129 601 5 N L=1.8e-07 W=1e-06 $X=299500 $Y=594385 $D=0
M4 602 134 5 5 N L=1.8e-07 W=1e-06 $X=300460 $Y=594385 $D=0
M5 123 132 602 5 N L=1.8e-07 W=1e-06 $X=301100 $Y=594385 $D=0
M6 603 132 123 5 N L=1.8e-07 W=1e-06 $X=301820 $Y=594385 $D=0
M7 5 134 603 5 N L=1.8e-07 W=1e-06 $X=302590 $Y=594385 $D=0
M8 79 472 5 5 N L=1.8e-07 W=1e-06 $X=325560 $Y=529975 $D=0
M9 5 472 79 5 N L=1.8e-07 W=1e-06 $X=326280 $Y=529975 $D=0
M10 79 472 5 5 N L=1.8e-07 W=1e-06 $X=327000 $Y=529975 $D=0
M11 5 472 79 5 N L=1.8e-07 W=1e-06 $X=327720 $Y=529975 $D=0
M12 472 121 5 5 N L=1.8e-07 W=5e-07 $X=328440 $Y=530475 $D=0
M13 5 8 472 5 N L=1.8e-07 W=5e-07 $X=329160 $Y=530475 $D=0
M14 472 8 5 5 N L=1.8e-07 W=5e-07 $X=329880 $Y=530475 $D=0
M15 5 121 472 5 N L=1.8e-07 W=5e-07 $X=330600 $Y=530475 $D=0
M16 123 129 455 1 P L=1.8e-07 W=1.37e-06 $X=297360 $Y=596245 $D=16
M17 455 127 123 1 P L=1.8e-07 W=1.37e-06 $X=298080 $Y=596245 $D=16
M18 123 127 455 1 P L=1.8e-07 W=1.37e-06 $X=298840 $Y=596245 $D=16
M19 455 129 123 1 P L=1.8e-07 W=1.37e-06 $X=299580 $Y=596245 $D=16
M20 1 134 455 1 P L=1.8e-07 W=1.37e-06 $X=300340 $Y=596245 $D=16
M21 455 132 1 1 P L=1.8e-07 W=1.37e-06 $X=301100 $Y=596245 $D=16
M22 1 132 455 1 P L=1.8e-07 W=1.37e-06 $X=301820 $Y=596245 $D=16
M23 455 134 1 1 P L=1.8e-07 W=1.37e-06 $X=302590 $Y=596245 $D=16
M24 79 472 1 1 P L=1.8e-07 W=1.37e-06 $X=325300 $Y=527745 $D=16
M25 1 472 79 1 P L=1.8e-07 W=1.37e-06 $X=326020 $Y=527745 $D=16
M26 79 472 1 1 P L=1.8e-07 W=1.37e-06 $X=326740 $Y=527745 $D=16
M27 1 472 79 1 P L=1.8e-07 W=1.37e-06 $X=327460 $Y=527745 $D=16
M28 604 121 1 1 P L=1.8e-07 W=1.37e-06 $X=328440 $Y=527745 $D=16
M29 472 8 604 1 P L=1.8e-07 W=1.37e-06 $X=329160 $Y=527745 $D=16
M30 605 8 472 1 P L=1.8e-07 W=1.37e-06 $X=329880 $Y=527745 $D=16
M31 1 121 605 1 P L=1.8e-07 W=1.37e-06 $X=330600 $Y=527745 $D=16
X215 1 5 DCAPBWP7T $T=156120 484280 0 0 $X=155830 $Y=484045
X216 1 5 DCAPBWP7T $T=165640 547000 1 0 $X=165350 $Y=542790
X217 1 5 DCAPBWP7T $T=177400 578360 0 0 $X=177110 $Y=578125
X218 1 5 DCAPBWP7T $T=185240 586200 0 0 $X=184950 $Y=585965
X219 1 5 DCAPBWP7T $T=188600 515640 1 0 $X=188310 $Y=511430
X220 1 5 DCAPBWP7T $T=195320 578360 0 0 $X=195030 $Y=578125
X221 1 5 DCAPBWP7T $T=195320 586200 0 0 $X=195030 $Y=585965
X222 1 5 DCAPBWP7T $T=220520 594040 0 0 $X=220230 $Y=593805
X223 1 5 DCAPBWP7T $T=226120 531320 0 0 $X=225830 $Y=531085
X224 1 5 DCAPBWP7T $T=237320 547000 1 0 $X=237030 $Y=542790
X225 1 5 DCAPBWP7T $T=237320 578360 1 0 $X=237030 $Y=574150
X226 1 5 DCAPBWP7T $T=237320 594040 0 0 $X=237030 $Y=593805
X227 1 5 DCAPBWP7T $T=251320 594040 1 0 $X=251030 $Y=589830
X228 1 5 DCAPBWP7T $T=264760 570520 0 0 $X=264470 $Y=570285
X229 1 5 DCAPBWP7T $T=267560 515640 0 0 $X=267270 $Y=515405
X230 1 5 DCAPBWP7T $T=279320 578360 0 0 $X=279030 $Y=578125
X231 1 5 DCAPBWP7T $T=279320 594040 1 0 $X=279030 $Y=589830
X232 1 5 DCAPBWP7T $T=282120 523480 1 0 $X=281830 $Y=519270
X233 1 5 DCAPBWP7T $T=291080 499960 0 0 $X=290790 $Y=499725
X234 1 5 DCAPBWP7T $T=293320 554840 0 0 $X=293030 $Y=554605
X235 1 5 DCAPBWP7T $T=293320 586200 1 0 $X=293030 $Y=581990
X236 1 5 DCAPBWP7T $T=306760 578360 1 0 $X=306470 $Y=574150
X237 1 5 DCAPBWP7T $T=309000 547000 0 0 $X=308710 $Y=546765
X238 1 5 DCAPBWP7T $T=321320 499960 0 0 $X=321030 $Y=499725
X239 1 5 DCAPBWP7T $T=321320 523480 0 0 $X=321030 $Y=523245
X240 1 5 DCAPBWP7T $T=321320 531320 1 0 $X=321030 $Y=527110
X241 1 5 DCAPBWP7T $T=324120 499960 0 0 $X=323830 $Y=499725
X242 1 5 DCAPBWP7T $T=324120 547000 0 0 $X=323830 $Y=546765
X243 1 5 DCAPBWP7T $T=334200 547000 0 0 $X=333910 $Y=546765
X244 1 5 DCAPBWP7T $T=335320 523480 1 0 $X=335030 $Y=519270
X245 1 5 DCAPBWP7T $T=338120 570520 1 0 $X=337830 $Y=566310
X246 1 5 DCAPBWP7T $T=339800 539160 0 0 $X=339510 $Y=538925
X247 1 5 DCAPBWP7T $T=347640 531320 0 0 $X=347350 $Y=531085
X248 1 5 DCAPBWP7T $T=354360 539160 0 0 $X=354070 $Y=538925
X249 1 5 DCAPBWP7T $T=363320 492120 1 0 $X=363030 $Y=487910
X250 1 5 DCAPBWP7T $T=363320 531320 1 0 $X=363030 $Y=527110
X251 1 5 DCAPBWP7T $T=363320 562680 0 0 $X=363030 $Y=562445
X252 1 5 DCAPBWP7T $T=363320 578360 0 0 $X=363030 $Y=578125
X253 1 5 DCAPBWP7T $T=366120 539160 0 0 $X=365830 $Y=538925
X254 1 5 DCAPBWP7T $T=372840 531320 1 0 $X=372550 $Y=527110
X255 1 5 DCAPBWP7T $T=381800 578360 0 0 $X=381510 $Y=578125
X256 1 5 DCAPBWP7T $T=390200 523480 0 0 $X=389910 $Y=523245
X257 1 5 DCAPBWP7T $T=405320 531320 1 0 $X=405030 $Y=527110
X258 1 5 DCAPBWP7T $T=405320 539160 0 0 $X=405030 $Y=538925
X259 1 5 DCAPBWP7T $T=405320 586200 0 0 $X=405030 $Y=585965
X260 1 5 DCAPBWP7T $T=405320 594040 1 0 $X=405030 $Y=589830
X261 1 5 DCAPBWP7T $T=405320 594040 0 0 $X=405030 $Y=593805
X262 1 5 DCAPBWP7T $T=412600 586200 1 0 $X=412310 $Y=581990
X263 1 5 DCAPBWP7T $T=421560 554840 0 0 $X=421270 $Y=554605
X264 1 5 DCAPBWP7T $T=427160 586200 1 0 $X=426870 $Y=581990
X265 1 5 DCAPBWP7T $T=431080 515640 0 0 $X=430790 $Y=515405
X266 1 5 DCAPBWP7T $T=439480 586200 0 0 $X=439190 $Y=585965
X267 1 5 DCAPBWP7T $T=439480 594040 0 0 $X=439190 $Y=593805
X268 1 5 DCAPBWP7T $T=447320 547000 0 0 $X=447030 $Y=546765
X269 5 1 DCAP8BWP7T $T=156120 578360 0 0 $X=155830 $Y=578125
X270 5 1 DCAP8BWP7T $T=156120 594040 1 0 $X=155830 $Y=589830
X271 5 1 DCAP8BWP7T $T=161160 547000 1 0 $X=160870 $Y=542790
X272 5 1 DCAP8BWP7T $T=174040 492120 1 0 $X=173750 $Y=487910
X273 5 1 DCAP8BWP7T $T=181320 578360 0 0 $X=181030 $Y=578125
X274 5 1 DCAP8BWP7T $T=182440 499960 0 0 $X=182150 $Y=499725
X275 5 1 DCAP8BWP7T $T=191400 492120 1 0 $X=191110 $Y=487910
X276 5 1 DCAP8BWP7T $T=191960 499960 0 0 $X=191670 $Y=499725
X277 5 1 DCAP8BWP7T $T=191960 523480 1 0 $X=191670 $Y=519270
X278 5 1 DCAP8BWP7T $T=191960 570520 1 0 $X=191670 $Y=566310
X279 5 1 DCAP8BWP7T $T=192520 562680 1 0 $X=192230 $Y=558470
X280 5 1 DCAP8BWP7T $T=216040 547000 0 0 $X=215750 $Y=546765
X281 5 1 DCAP8BWP7T $T=216040 562680 0 0 $X=215750 $Y=562445
X282 5 1 DCAP8BWP7T $T=216040 594040 0 0 $X=215750 $Y=593805
X283 5 1 DCAP8BWP7T $T=232840 578360 1 0 $X=232550 $Y=574150
X284 5 1 DCAP8BWP7T $T=232840 594040 0 0 $X=232550 $Y=593805
X285 5 1 DCAP8BWP7T $T=233400 499960 0 0 $X=233110 $Y=499725
X286 5 1 DCAP8BWP7T $T=233960 507800 1 0 $X=233670 $Y=503590
X287 5 1 DCAP8BWP7T $T=234520 515640 1 0 $X=234230 $Y=511430
X288 5 1 DCAP8BWP7T $T=234520 562680 0 0 $X=234230 $Y=562445
X289 5 1 DCAP8BWP7T $T=275960 531320 1 0 $X=275670 $Y=527110
X290 5 1 DCAP8BWP7T $T=275960 547000 0 0 $X=275670 $Y=546765
X291 5 1 DCAP8BWP7T $T=275960 586200 1 0 $X=275670 $Y=581990
X292 5 1 DCAP8BWP7T $T=275960 586200 0 0 $X=275670 $Y=585965
X293 5 1 DCAP8BWP7T $T=276520 499960 1 0 $X=276230 $Y=495750
X294 5 1 DCAP8BWP7T $T=285480 515640 0 0 $X=285190 $Y=515405
X295 5 1 DCAP8BWP7T $T=289960 507800 1 0 $X=289670 $Y=503590
X296 5 1 DCAP8BWP7T $T=303400 594040 0 0 $X=303110 $Y=593805
X297 5 1 DCAP8BWP7T $T=307880 554840 0 0 $X=307590 $Y=554605
X298 5 1 DCAP8BWP7T $T=308440 492120 0 0 $X=308150 $Y=491885
X299 5 1 DCAP8BWP7T $T=318520 515640 0 0 $X=318230 $Y=515405
X300 5 1 DCAP8BWP7T $T=324120 507800 0 0 $X=323830 $Y=507565
X301 5 1 DCAP8BWP7T $T=324120 586200 0 0 $X=323830 $Y=585965
X302 5 1 DCAP8BWP7T $T=335320 570520 0 0 $X=335030 $Y=570285
X303 5 1 DCAP8BWP7T $T=335320 586200 1 0 $X=335030 $Y=581990
X304 5 1 DCAP8BWP7T $T=343160 531320 0 0 $X=342870 $Y=531085
X305 5 1 DCAP8BWP7T $T=359960 492120 0 0 $X=359670 $Y=491885
X306 5 1 DCAP8BWP7T $T=359960 578360 1 0 $X=359670 $Y=574150
X307 5 1 DCAP8BWP7T $T=359960 594040 0 0 $X=359670 $Y=593805
X308 5 1 DCAP8BWP7T $T=366120 499960 1 0 $X=365830 $Y=495750
X309 5 1 DCAP8BWP7T $T=377880 507800 1 0 $X=377590 $Y=503590
X310 5 1 DCAP8BWP7T $T=384040 547000 0 0 $X=383750 $Y=546765
X311 5 1 DCAP8BWP7T $T=389640 507800 1 0 $X=389350 $Y=503590
X312 5 1 DCAP8BWP7T $T=401960 507800 0 0 $X=401670 $Y=507565
X313 5 1 DCAP8BWP7T $T=401960 562680 0 0 $X=401670 $Y=562445
X314 5 1 DCAP8BWP7T $T=401960 570520 0 0 $X=401670 $Y=570285
X315 5 1 DCAP8BWP7T $T=401960 578360 1 0 $X=401670 $Y=574150
X316 5 1 DCAP8BWP7T $T=408120 531320 0 0 $X=407830 $Y=531085
X317 5 1 DCAP8BWP7T $T=408120 586200 1 0 $X=407830 $Y=581990
X318 5 1 DCAP8BWP7T $T=443400 515640 0 0 $X=443110 $Y=515405
X319 5 1 DCAP8BWP7T $T=443400 531320 0 0 $X=443110 $Y=531085
X320 5 1 DCAP8BWP7T $T=444520 484280 0 0 $X=444230 $Y=484045
X321 5 1 DCAP8BWP7T $T=444520 499960 0 0 $X=444230 $Y=499725
X322 5 1 DCAP8BWP7T $T=444520 554840 0 0 $X=444230 $Y=554605
X323 5 1 DCAP8BWP7T $T=444520 578360 1 0 $X=444230 $Y=574150
X324 5 1 DCAP8BWP7T $T=444520 578360 0 0 $X=444230 $Y=578125
X325 5 1 DCAP8BWP7T $T=444520 586200 0 0 $X=444230 $Y=585965
X326 5 1 DCAP4BWP7T $T=165080 507800 0 0 $X=164790 $Y=507565
X327 5 1 DCAP4BWP7T $T=169000 484280 0 0 $X=168710 $Y=484045
X328 5 1 DCAP4BWP7T $T=183000 586200 0 0 $X=182710 $Y=585965
X329 5 1 DCAP4BWP7T $T=188040 570520 1 0 $X=187750 $Y=566310
X330 5 1 DCAP4BWP7T $T=193080 578360 0 0 $X=192790 $Y=578125
X331 5 1 DCAP4BWP7T $T=194200 492120 0 0 $X=193910 $Y=491885
X332 5 1 DCAP4BWP7T $T=194760 484280 0 0 $X=194470 $Y=484045
X333 5 1 DCAP4BWP7T $T=194760 515640 0 0 $X=194470 $Y=515405
X334 5 1 DCAP4BWP7T $T=236200 562680 1 0 $X=235910 $Y=558470
X335 5 1 DCAP4BWP7T $T=236200 570520 1 0 $X=235910 $Y=566310
X336 5 1 DCAP4BWP7T $T=249080 570520 1 0 $X=248790 $Y=566310
X337 5 1 DCAP4BWP7T $T=253560 515640 1 0 $X=253270 $Y=511430
X338 5 1 DCAP4BWP7T $T=253560 578360 0 0 $X=253270 $Y=578125
X339 5 1 DCAP4BWP7T $T=267000 507800 0 0 $X=266710 $Y=507565
X340 5 1 DCAP4BWP7T $T=291080 554840 0 0 $X=290790 $Y=554605
X341 5 1 DCAP4BWP7T $T=291080 586200 1 0 $X=290790 $Y=581990
X342 5 1 DCAP4BWP7T $T=296120 570520 1 0 $X=295830 $Y=566310
X343 5 1 DCAP4BWP7T $T=302280 515640 1 0 $X=301990 $Y=511430
X344 5 1 DCAP4BWP7T $T=319080 523480 0 0 $X=318790 $Y=523245
X345 5 1 DCAP4BWP7T $T=319080 531320 1 0 $X=318790 $Y=527110
X346 5 1 DCAP4BWP7T $T=320200 531320 0 0 $X=319910 $Y=531085
X347 5 1 DCAP4BWP7T $T=320200 547000 1 0 $X=319910 $Y=542790
X348 5 1 DCAP4BWP7T $T=333080 523480 1 0 $X=332790 $Y=519270
X349 5 1 DCAP4BWP7T $T=335880 570520 1 0 $X=335590 $Y=566310
X350 5 1 DCAP4BWP7T $T=347640 523480 1 0 $X=347350 $Y=519270
X351 5 1 DCAP4BWP7T $T=361080 492120 1 0 $X=360790 $Y=487910
X352 5 1 DCAP4BWP7T $T=361080 531320 1 0 $X=360790 $Y=527110
X353 5 1 DCAP4BWP7T $T=362200 586200 0 0 $X=361910 $Y=585965
X354 5 1 DCAP4BWP7T $T=366120 507800 1 0 $X=365830 $Y=503590
X355 5 1 DCAP4BWP7T $T=366120 570520 1 0 $X=365830 $Y=566310
X356 5 1 DCAP4BWP7T $T=370040 586200 0 0 $X=369750 $Y=585965
X357 5 1 DCAP4BWP7T $T=387960 523480 0 0 $X=387670 $Y=523245
X358 5 1 DCAP4BWP7T $T=403080 586200 0 0 $X=402790 $Y=585965
X359 5 1 DCAP4BWP7T $T=404200 515640 1 0 $X=403910 $Y=511430
X360 5 1 DCAP4BWP7T $T=404760 499960 0 0 $X=404470 $Y=499725
X361 5 1 DCAP4BWP7T $T=404760 515640 0 0 $X=404470 $Y=515405
X362 5 1 DCAP4BWP7T $T=417080 492120 0 0 $X=416790 $Y=491885
X363 5 1 DCAP4BWP7T $T=437240 594040 0 0 $X=436950 $Y=593805
X364 5 1 DCAP4BWP7T $T=446760 492120 0 0 $X=446470 $Y=491885
X365 5 1 ICV_40 $T=174040 531320 1 0 $X=173750 $Y=527110
X366 5 1 ICV_40 $T=177400 578360 1 0 $X=177110 $Y=574150
X367 5 1 ICV_40 $T=183000 562680 1 0 $X=182710 $Y=558470
X368 5 1 ICV_40 $T=188600 586200 0 0 $X=188310 $Y=585965
X369 5 1 ICV_40 $T=189160 539160 1 0 $X=188870 $Y=534950
X370 5 1 ICV_40 $T=189720 547000 1 0 $X=189430 $Y=542790
X371 5 1 ICV_40 $T=189720 586200 1 0 $X=189430 $Y=581990
X372 5 1 ICV_40 $T=189720 594040 1 0 $X=189430 $Y=589830
X373 5 1 ICV_40 $T=190280 539160 0 0 $X=189990 $Y=538925
X374 5 1 ICV_40 $T=190280 562680 0 0 $X=189990 $Y=562445
X375 5 1 ICV_40 $T=198120 515640 0 0 $X=197830 $Y=515405
X376 5 1 ICV_40 $T=198120 578360 1 0 $X=197830 $Y=574150
X377 5 1 ICV_40 $T=207080 499960 0 0 $X=206790 $Y=499725
X378 5 1 ICV_40 $T=223320 507800 1 0 $X=223030 $Y=503590
X379 5 1 ICV_40 $T=230600 547000 1 0 $X=230310 $Y=542790
X380 5 1 ICV_40 $T=231160 554840 0 0 $X=230870 $Y=554605
X381 5 1 ICV_40 $T=231720 523480 0 0 $X=231430 $Y=523245
X382 5 1 ICV_40 $T=232280 515640 0 0 $X=231990 $Y=515405
X383 5 1 ICV_40 $T=232280 531320 1 0 $X=231990 $Y=527110
X384 5 1 ICV_40 $T=232280 539160 1 0 $X=231990 $Y=534950
X385 5 1 ICV_40 $T=258040 570520 0 0 $X=257750 $Y=570285
X386 5 1 ICV_40 $T=258040 594040 0 0 $X=257750 $Y=593805
X387 5 1 ICV_40 $T=272600 578360 0 0 $X=272310 $Y=578125
X388 5 1 ICV_40 $T=272600 594040 1 0 $X=272310 $Y=589830
X389 5 1 ICV_40 $T=273160 499960 0 0 $X=272870 $Y=499725
X390 5 1 ICV_40 $T=273720 539160 1 0 $X=273430 $Y=534950
X391 5 1 ICV_40 $T=273720 570520 0 0 $X=273430 $Y=570285
X392 5 1 ICV_40 $T=282120 515640 1 0 $X=281830 $Y=511430
X393 5 1 ICV_40 $T=291080 562680 0 0 $X=290790 $Y=562445
X394 5 1 ICV_40 $T=298920 507800 1 0 $X=298630 $Y=503590
X395 5 1 ICV_40 $T=300040 539160 1 0 $X=299750 $Y=534950
X396 5 1 ICV_40 $T=300040 578360 0 0 $X=299750 $Y=578125
X397 5 1 ICV_40 $T=300040 594040 1 0 $X=299750 $Y=589830
X398 5 1 ICV_40 $T=305080 570520 1 0 $X=304790 $Y=566310
X399 5 1 ICV_40 $T=308440 515640 0 0 $X=308150 $Y=515405
X400 5 1 ICV_40 $T=314600 499960 0 0 $X=314310 $Y=499725
X401 5 1 ICV_40 $T=315720 515640 1 0 $X=315430 $Y=511430
X402 5 1 ICV_40 $T=324120 492120 0 0 $X=323830 $Y=491885
X403 5 1 ICV_40 $T=324120 531320 0 0 $X=323830 $Y=531085
X404 5 1 ICV_40 $T=324120 570520 1 0 $X=323830 $Y=566310
X405 5 1 ICV_40 $T=330280 507800 0 0 $X=329990 $Y=507565
X406 5 1 ICV_40 $T=333080 539160 0 0 $X=332790 $Y=538925
X407 5 1 ICV_40 $T=340360 531320 1 0 $X=340070 $Y=527110
X408 5 1 ICV_40 $T=342040 515640 1 0 $X=341750 $Y=511430
X409 5 1 ICV_40 $T=350440 578360 1 0 $X=350150 $Y=574150
X410 5 1 ICV_40 $T=351000 515640 1 0 $X=350710 $Y=511430
X411 5 1 ICV_40 $T=357720 515640 0 0 $X=357430 $Y=515405
X412 5 1 ICV_40 $T=357720 594040 1 0 $X=357430 $Y=589830
X413 5 1 ICV_40 $T=358280 499960 1 0 $X=357990 $Y=495750
X414 5 1 ICV_40 $T=358280 570520 0 0 $X=357990 $Y=570285
X415 5 1 ICV_40 $T=366120 492120 1 0 $X=365830 $Y=487910
X416 5 1 ICV_40 $T=366120 531320 1 0 $X=365830 $Y=527110
X417 5 1 ICV_40 $T=375080 499960 0 0 $X=374790 $Y=499725
X418 5 1 ICV_40 $T=377880 594040 1 0 $X=377590 $Y=589830
X419 5 1 ICV_40 $T=398600 539160 0 0 $X=398310 $Y=538925
X420 5 1 ICV_40 $T=398600 594040 1 0 $X=398310 $Y=589830
X421 5 1 ICV_40 $T=424360 515640 0 0 $X=424070 $Y=515405
X422 5 1 ICV_40 $T=440600 547000 0 0 $X=440310 $Y=546765
X423 5 1 ICV_40 $T=441160 515640 1 0 $X=440870 $Y=511430
X424 5 1 ICV_40 $T=441160 531320 1 0 $X=440870 $Y=527110
X425 5 1 ICV_40 $T=441720 507800 1 0 $X=441430 $Y=503590
X426 5 1 ICV_40 $T=441720 554840 1 0 $X=441430 $Y=550630
X427 5 1 ICV_40 $T=441720 586200 1 0 $X=441430 $Y=581990
X428 5 1 ICV_40 $T=442280 499960 1 0 $X=441990 $Y=495750
X429 5 1 ICV_40 $T=442280 547000 1 0 $X=441990 $Y=542790
X430 284 1 281 8 5 NR2D1BWP7T $T=158360 515640 0 180 $X=155830 $Y=511430
X431 10 1 290 8 5 NR2D1BWP7T $T=158920 547000 1 0 $X=158630 $Y=542790
X432 15 1 291 12 5 NR2D1BWP7T $T=161720 586200 0 180 $X=159190 $Y=581990
X433 10 1 292 17 5 NR2D1BWP7T $T=159480 594040 0 0 $X=159190 $Y=593805
X434 20 1 289 8 5 NR2D1BWP7T $T=163960 578360 1 180 $X=161430 $Y=578125
X435 22 1 296 20 5 NR2D1BWP7T $T=163960 594040 1 180 $X=161430 $Y=593805
X436 12 1 298 8 5 NR2D1BWP7T $T=164520 562680 0 0 $X=164230 $Y=562445
X437 25 1 297 8 5 NR2D1BWP7T $T=167880 515640 1 180 $X=165350 $Y=515405
X438 33 1 301 8 5 NR2D1BWP7T $T=172360 562680 1 180 $X=169830 $Y=562445
X439 35 1 302 8 5 NR2D1BWP7T $T=175160 578360 0 180 $X=172630 $Y=574150
X440 307 1 287 8 5 NR2D1BWP7T $T=177400 578360 0 180 $X=174870 $Y=574150
X441 315 1 308 8 5 NR2D1BWP7T $T=179080 570520 0 180 $X=176550 $Y=566310
X442 41 1 288 8 5 NR2D1BWP7T $T=180760 523480 0 180 $X=178230 $Y=519270
X443 318 1 309 8 5 NR2D1BWP7T $T=180760 570520 1 180 $X=178230 $Y=570285
X444 284 1 313 310 5 NR2D1BWP7T $T=181320 515640 0 180 $X=178790 $Y=511430
X445 307 1 314 316 5 NR2D1BWP7T $T=179080 539160 0 0 $X=178790 $Y=538925
X446 42 1 312 307 5 NR2D1BWP7T $T=181320 578360 1 180 $X=178790 $Y=578125
X447 316 1 40 8 5 NR2D1BWP7T $T=181880 507800 0 180 $X=179350 $Y=503590
X448 42 1 321 284 5 NR2D1BWP7T $T=184120 507800 0 180 $X=181590 $Y=503590
X449 320 1 322 307 5 NR2D1BWP7T $T=181880 570520 1 0 $X=181590 $Y=566310
X450 284 1 323 316 5 NR2D1BWP7T $T=182440 515640 1 0 $X=182150 $Y=511430
X451 318 1 325 332 5 NR2D1BWP7T $T=184680 578360 1 0 $X=184390 $Y=574150
X452 326 1 329 336 5 NR2D1BWP7T $T=185800 554840 1 0 $X=185510 $Y=550630
X453 326 1 330 332 5 NR2D1BWP7T $T=185800 570520 1 0 $X=185510 $Y=566310
X454 318 1 331 320 5 NR2D1BWP7T $T=189160 539160 0 180 $X=186630 $Y=534950
X455 326 1 337 8 5 NR2D1BWP7T $T=189720 547000 0 180 $X=187190 $Y=542790
X456 326 1 338 310 5 NR2D1BWP7T $T=190280 507800 0 180 $X=187750 $Y=503590
X457 318 1 341 310 5 NR2D1BWP7T $T=192520 507800 0 180 $X=189990 $Y=503590
X458 336 1 55 8 5 NR2D1BWP7T $T=192520 515640 0 180 $X=189990 $Y=511430
X459 42 1 343 35 5 NR2D1BWP7T $T=190280 570520 0 0 $X=189990 $Y=570285
X460 315 1 345 332 5 NR2D1BWP7T $T=198680 531320 0 0 $X=198390 $Y=531085
X461 315 1 351 310 5 NR2D1BWP7T $T=204840 523480 1 0 $X=204550 $Y=519270
X462 310 1 62 8 5 NR2D1BWP7T $T=213240 499960 0 180 $X=210710 $Y=495750
X463 35 1 74 316 5 NR2D1BWP7T $T=218280 570520 1 180 $X=215750 $Y=570285
X464 315 1 363 320 5 NR2D1BWP7T $T=226120 539160 1 0 $X=225830 $Y=534950
X465 320 1 377 284 5 NR2D1BWP7T $T=230040 531320 1 180 $X=227510 $Y=531085
X466 315 1 383 316 5 NR2D1BWP7T $T=229480 523480 0 0 $X=229190 $Y=523245
X467 326 1 382 320 5 NR2D1BWP7T $T=232280 515640 0 180 $X=229750 $Y=511430
X468 318 1 385 316 5 NR2D1BWP7T $T=231160 499960 0 0 $X=230870 $Y=499725
X469 42 1 387 315 5 NR2D1BWP7T $T=234520 515640 0 180 $X=231990 $Y=511430
X470 336 1 434 318 5 NR2D1BWP7T $T=274280 515640 1 0 $X=273990 $Y=511430
X471 326 1 438 42 5 NR2D1BWP7T $T=283240 515640 0 0 $X=282950 $Y=515405
X472 117 1 116 115 5 NR2D1BWP7T $T=287720 594040 1 180 $X=285190 $Y=593805
X473 42 1 417 318 5 NR2D1BWP7T $T=306760 515640 0 180 $X=304230 $Y=511430
X474 156 1 457 8 5 NR2D1BWP7T $T=329160 492120 1 0 $X=328870 $Y=487910
X475 168 1 475 8 5 NR2D1BWP7T $T=337560 515640 1 180 $X=335030 $Y=515405
X476 162 1 483 164 5 NR2D1BWP7T $T=335880 547000 0 0 $X=335590 $Y=546765
X477 165 1 465 115 5 NR2D1BWP7T $T=340360 586200 1 180 $X=337830 $Y=585965
X478 166 1 488 168 5 NR2D1BWP7T $T=339800 570520 1 0 $X=339510 $Y=566310
X479 167 1 456 115 5 NR2D1BWP7T $T=342040 586200 0 180 $X=339510 $Y=581990
X480 170 1 169 8 5 NR2D1BWP7T $T=343160 492120 0 180 $X=340630 $Y=487910
X481 162 1 484 172 5 NR2D1BWP7T $T=342600 570520 0 0 $X=342310 $Y=570285
X482 162 1 492 8 5 NR2D1BWP7T $T=348760 515640 1 180 $X=346230 $Y=515405
X483 172 1 496 168 5 NR2D1BWP7T $T=348760 578360 1 180 $X=346230 $Y=578125
X484 172 1 498 173 5 NR2D1BWP7T $T=347080 570520 0 0 $X=346790 $Y=570285
X485 166 1 494 170 5 NR2D1BWP7T $T=349880 562680 1 180 $X=347350 $Y=562445
X486 176 1 489 173 5 NR2D1BWP7T $T=350440 570520 0 180 $X=347910 $Y=566310
X487 173 1 491 8 5 NR2D1BWP7T $T=351000 515640 0 180 $X=348470 $Y=511430
X488 166 1 178 115 5 NR2D1BWP7T $T=352680 586200 0 180 $X=350150 $Y=581990
X489 181 1 179 8 5 NR2D1BWP7T $T=353240 507800 0 180 $X=350710 $Y=503590
X490 183 1 476 8 5 NR2D1BWP7T $T=356040 507800 0 180 $X=353510 $Y=503590
X491 166 1 517 162 5 NR2D1BWP7T $T=368920 594040 0 180 $X=366390 $Y=589830
X492 162 1 468 176 5 NR2D1BWP7T $T=367240 578360 0 0 $X=366950 $Y=578125
X493 176 1 497 168 5 NR2D1BWP7T $T=368920 578360 1 0 $X=368630 $Y=574150
X494 166 1 520 183 5 NR2D1BWP7T $T=372840 578360 1 180 $X=370310 $Y=578125
X495 193 1 519 8 5 NR2D1BWP7T $T=373400 492120 1 180 $X=370870 $Y=491885
X496 195 1 525 202 5 NR2D1BWP7T $T=372840 492120 1 0 $X=372550 $Y=487910
X497 164 1 526 173 5 NR2D1BWP7T $T=373400 570520 1 0 $X=373110 $Y=566310
X498 172 1 534 170 5 NR2D1BWP7T $T=382360 578360 0 180 $X=379830 $Y=574150
X499 176 1 535 183 5 NR2D1BWP7T $T=385720 578360 1 180 $X=383190 $Y=578125
X500 181 1 555 176 5 NR2D1BWP7T $T=401960 562680 1 180 $X=399430 $Y=562445
X501 195 1 550 8 5 NR2D1BWP7T $T=417640 515640 0 180 $X=415110 $Y=511430
X502 230 1 570 8 5 NR2D1BWP7T $T=424360 499960 0 180 $X=421830 $Y=495750
X503 176 1 528 170 5 NR2D1BWP7T $T=424920 578360 1 180 $X=422390 $Y=578125
X504 172 1 553 183 5 NR2D1BWP7T $T=427160 594040 0 0 $X=426870 $Y=593805
X505 244 1 545 8 5 NR2D1BWP7T $T=434440 531320 0 180 $X=431910 $Y=527110
X506 267 1 262 260 5 NR2D1BWP7T $T=444520 554840 1 180 $X=441990 $Y=554605
X507 268 1 254 260 5 NR2D1BWP7T $T=444520 578360 0 180 $X=441990 $Y=574150
X508 1 5 DCAP64BWP7T $T=158360 492120 0 0 $X=158070 $Y=491885
X509 1 5 DCAP64BWP7T $T=369480 594040 0 0 $X=369190 $Y=593805
X510 1 5 DCAP64BWP7T $T=408120 492120 1 0 $X=407830 $Y=487910
X511 1 5 DCAP64BWP7T $T=408120 507800 0 0 $X=407830 $Y=507565
X512 1 5 DCAP64BWP7T $T=408120 523480 0 0 $X=407830 $Y=523245
X513 1 5 DCAP64BWP7T $T=408120 539160 1 0 $X=407830 $Y=534950
X514 1 5 DCAP64BWP7T $T=408120 539160 0 0 $X=407830 $Y=538925
X515 1 5 DCAP64BWP7T $T=408120 562680 0 0 $X=407830 $Y=562445
X516 1 5 DCAP64BWP7T $T=408120 594040 1 0 $X=407830 $Y=589830
X564 5 1 ICV_47 $T=156120 523480 0 0 $X=155830 $Y=523245
X565 5 1 ICV_47 $T=156120 547000 0 0 $X=155830 $Y=546765
X566 5 1 ICV_47 $T=198120 492120 0 0 $X=197830 $Y=491885
X567 5 1 ICV_47 $T=198120 507800 0 0 $X=197830 $Y=507565
X568 5 1 ICV_47 $T=198120 578360 0 0 $X=197830 $Y=578125
X569 5 1 ICV_47 $T=198120 594040 1 0 $X=197830 $Y=589830
X570 5 1 ICV_47 $T=240120 492120 1 0 $X=239830 $Y=487910
X571 5 1 ICV_47 $T=240120 492120 0 0 $X=239830 $Y=491885
X572 5 1 ICV_47 $T=240120 507800 1 0 $X=239830 $Y=503590
X573 5 1 ICV_47 $T=240120 523480 1 0 $X=239830 $Y=519270
X574 5 1 ICV_47 $T=240120 531320 0 0 $X=239830 $Y=531085
X575 5 1 ICV_47 $T=240120 547000 1 0 $X=239830 $Y=542790
X576 5 1 ICV_47 $T=240120 562680 1 0 $X=239830 $Y=558470
X577 5 1 ICV_47 $T=282120 484280 0 0 $X=281830 $Y=484045
X578 5 1 ICV_47 $T=282120 507800 0 0 $X=281830 $Y=507565
X579 5 1 ICV_47 $T=324120 484280 0 0 $X=323830 $Y=484045
X580 5 1 ICV_47 $T=324120 523480 0 0 $X=323830 $Y=523245
X581 5 1 ICV_47 $T=324120 539160 1 0 $X=323830 $Y=534950
X582 5 1 ICV_47 $T=324120 554840 1 0 $X=323830 $Y=550630
X583 5 1 ICV_47 $T=324120 562680 1 0 $X=323830 $Y=558470
X584 5 1 ICV_47 $T=366120 484280 0 0 $X=365830 $Y=484045
X585 5 1 ICV_47 $T=366120 523480 1 0 $X=365830 $Y=519270
X586 5 1 ICV_47 $T=366120 531320 0 0 $X=365830 $Y=531085
X587 5 1 ICV_47 $T=366120 547000 1 0 $X=365830 $Y=542790
X588 5 1 ICV_47 $T=366120 554840 0 0 $X=365830 $Y=554605
X589 5 1 ICV_47 $T=366120 586200 1 0 $X=365830 $Y=581990
X590 1 5 DCAP32BWP7T $T=158360 515640 1 0 $X=158070 $Y=511430
X591 1 5 DCAP32BWP7T $T=167880 515640 0 0 $X=167590 $Y=515405
X592 1 5 DCAP32BWP7T $T=174600 507800 0 0 $X=174310 $Y=507565
X593 1 5 DCAP32BWP7T $T=175720 499960 1 0 $X=175430 $Y=495750
X594 1 5 DCAP32BWP7T $T=176840 484280 0 0 $X=176550 $Y=484045
X595 1 5 DCAP32BWP7T $T=198120 515640 1 0 $X=197830 $Y=511430
X596 1 5 DCAP32BWP7T $T=198120 547000 0 0 $X=197830 $Y=546765
X597 1 5 DCAP32BWP7T $T=198120 570520 0 0 $X=197830 $Y=570285
X598 1 5 DCAP32BWP7T $T=209320 562680 1 0 $X=209030 $Y=558470
X599 1 5 DCAP32BWP7T $T=221080 484280 0 0 $X=220790 $Y=484045
X600 1 5 DCAP32BWP7T $T=240120 507800 0 0 $X=239830 $Y=507565
X601 1 5 DCAP32BWP7T $T=253560 562680 0 0 $X=253270 $Y=562445
X602 1 5 DCAP32BWP7T $T=282120 539160 1 0 $X=281830 $Y=534950
X603 1 5 DCAP32BWP7T $T=282120 547000 0 0 $X=281830 $Y=546765
X604 1 5 DCAP32BWP7T $T=287720 531320 0 0 $X=287430 $Y=531085
X605 1 5 DCAP32BWP7T $T=291080 499960 1 0 $X=290790 $Y=495750
X606 1 5 DCAP32BWP7T $T=295560 562680 1 0 $X=295270 $Y=558470
X607 1 5 DCAP32BWP7T $T=301160 531320 1 0 $X=300870 $Y=527110
X608 1 5 DCAP32BWP7T $T=301720 586200 0 0 $X=301430 $Y=585965
X609 1 5 DCAP32BWP7T $T=324120 507800 1 0 $X=323830 $Y=503590
X610 1 5 DCAP32BWP7T $T=324120 515640 1 0 $X=323830 $Y=511430
X611 1 5 DCAP32BWP7T $T=324120 562680 0 0 $X=323830 $Y=562445
X612 1 5 DCAP32BWP7T $T=324120 594040 1 0 $X=323830 $Y=589830
X613 1 5 DCAP32BWP7T $T=336440 499960 0 0 $X=336150 $Y=499725
X614 1 5 DCAP32BWP7T $T=344280 586200 0 0 $X=343990 $Y=585965
X615 1 5 DCAP32BWP7T $T=366120 562680 1 0 $X=365830 $Y=558470
X616 1 5 DCAP32BWP7T $T=375080 499960 1 0 $X=374790 $Y=495750
X617 1 5 DCAP32BWP7T $T=375640 570520 1 0 $X=375350 $Y=566310
X618 1 5 DCAP32BWP7T $T=380680 539160 0 0 $X=380390 $Y=538925
X619 1 5 DCAP32BWP7T $T=385160 586200 0 0 $X=384870 $Y=585965
X620 1 5 DCAP32BWP7T $T=385720 578360 0 0 $X=385430 $Y=578125
X621 1 5 DCAP32BWP7T $T=386840 499960 0 0 $X=386550 $Y=499725
X622 1 5 DCAP32BWP7T $T=408120 547000 0 0 $X=407830 $Y=546765
X623 1 5 DCAP32BWP7T $T=408120 578360 1 0 $X=407830 $Y=574150
X624 1 5 DCAP32BWP7T $T=417640 515640 1 0 $X=417350 $Y=511430
X625 1 5 DCAP32BWP7T $T=421560 562680 1 0 $X=421270 $Y=558470
X626 1 5 DCAP32BWP7T $T=421560 570520 0 0 $X=421270 $Y=570285
X627 1 5 DCAP32BWP7T $T=421560 586200 0 0 $X=421270 $Y=585965
X628 1 5 DCAP32BWP7T $T=424360 499960 1 0 $X=424070 $Y=495750
X629 291 292 296 311 1 5 317 FA1D0BWP7T $T=167880 594040 1 0 $X=167590 $Y=589830
X630 37 43 295 53 1 5 340 FA1D0BWP7T $T=178520 492120 1 0 $X=178230 $Y=487910
X631 306 304 348 68 1 5 357 FA1D0BWP7T $T=198680 492120 1 0 $X=198390 $Y=487910
X632 328 311 333 347 1 5 360 FA1D0BWP7T $T=198680 547000 1 0 $X=198390 $Y=542790
X633 324 57 64 359 1 5 69 FA1D0BWP7T $T=198680 586200 0 0 $X=198390 $Y=585965
X634 63 317 359 368 1 5 361 FA1D0BWP7T $T=209320 554840 0 0 $X=209030 $Y=554605
X635 312 363 330 370 1 5 371 FA1D0BWP7T $T=210440 531320 1 0 $X=210150 $Y=527110
X636 362 354 341 372 1 5 374 FA1D0BWP7T $T=213240 515640 0 0 $X=212950 $Y=515405
X637 331 321 338 373 1 5 376 FA1D0BWP7T $T=214920 499960 0 0 $X=214630 $Y=499725
X638 356 373 378 87 1 5 388 FA1D0BWP7T $T=221640 492120 1 0 $X=221350 $Y=487910
X639 343 325 329 386 1 5 393 FA1D0BWP7T $T=221640 547000 0 0 $X=221350 $Y=546765
X640 360 352 368 355 1 5 364 FA1D0BWP7T $T=221640 562680 0 0 $X=221350 $Y=562445
X641 370 376 372 397 1 5 96 FA1D0BWP7T $T=240680 499960 1 0 $X=240390 $Y=495750
X642 389 391 374 93 1 5 401 FA1D0BWP7T $T=240680 515640 1 0 $X=240390 $Y=511430
X643 353 351 377 391 1 5 403 FA1D0BWP7T $T=240680 523480 0 0 $X=240390 $Y=523245
X644 339 386 371 389 1 5 400 FA1D0BWP7T $T=240680 539160 1 0 $X=240390 $Y=534950
X645 313 322 345 394 1 5 402 FA1D0BWP7T $T=240680 554840 1 0 $X=240390 $Y=550630
X646 88 375 335 398 1 5 365 FA1D0BWP7T $T=240680 562680 0 0 $X=240390 $Y=562445
X647 390 90 92 381 1 5 94 FA1D0BWP7T $T=240680 578360 0 0 $X=240390 $Y=578125
X648 394 403 408 404 1 5 414 FA1D0BWP7T $T=250200 531320 1 0 $X=249910 $Y=527110
X649 395 404 400 412 1 5 410 FA1D0BWP7T $T=250760 539160 0 0 $X=250470 $Y=538925
X650 393 334 99 395 1 5 415 FA1D0BWP7T $T=250760 554840 0 0 $X=250470 $Y=554605
X651 396 385 387 413 1 5 101 FA1D0BWP7T $T=251320 499960 0 0 $X=251030 $Y=499725
X652 388 98 397 102 1 5 103 FA1D0BWP7T $T=253000 484280 0 0 $X=252710 $Y=484045
X653 100 412 401 432 1 5 435 FA1D0BWP7T $T=263080 531320 1 0 $X=262790 $Y=527110
X654 418 423 431 108 1 5 433 FA1D0BWP7T $T=263640 499960 1 0 $X=263350 $Y=495750
X655 434 428 422 408 1 5 399 FA1D0BWP7T $T=276520 554840 1 180 $X=263350 $Y=554605
X656 495 489 484 480 1 5 478 FA1D0BWP7T $T=347640 554840 1 180 $X=334470 $Y=554605
X657 487 481 482 499 1 5 500 FA1D0BWP7T $T=341480 539160 0 0 $X=341190 $Y=538925
X658 497 483 494 510 1 5 515 FA1D0BWP7T $T=347640 554840 0 0 $X=347350 $Y=554605
X659 513 521 528 530 1 5 531 FA1D0BWP7T $T=366680 554840 1 0 $X=366390 $Y=550630
X660 516 510 514 508 1 5 533 FA1D0BWP7T $T=367800 539160 0 0 $X=367510 $Y=538925
X661 194 496 520 532 1 5 537 FA1D0BWP7T $T=372280 586200 0 0 $X=371990 $Y=585965
X662 199 203 539 540 1 5 541 FA1D0BWP7T $T=376760 492120 0 0 $X=376470 $Y=491885
X663 532 515 530 543 1 5 546 FA1D0BWP7T $T=379560 554840 1 0 $X=379270 $Y=550630
X664 533 503 543 544 1 5 547 FA1D0BWP7T $T=380120 539160 1 0 $X=379830 $Y=534950
X665 527 534 212 548 1 5 549 FA1D0BWP7T $T=381240 562680 0 0 $X=380950 $Y=562445
X666 209 535 215 551 1 5 216 FA1D0BWP7T $T=385720 594040 1 0 $X=385430 $Y=589830
X667 210 213 553 554 1 5 559 FA1D0BWP7T $T=389080 578360 1 0 $X=388790 $Y=574150
X668 211 214 217 539 1 5 562 FA1D0BWP7T $T=389640 492120 0 0 $X=389350 $Y=491885
X669 542 548 531 557 1 5 563 FA1D0BWP7T $T=389640 547000 0 0 $X=389350 $Y=546765
X670 221 525 224 578 1 5 228 FA1D0BWP7T $T=408680 484280 0 0 $X=408390 $Y=484045
X671 578 574 223 568 1 5 564 FA1D0BWP7T $T=421560 499960 1 180 $X=408390 $Y=499725
X672 567 571 563 579 1 5 582 FA1D0BWP7T $T=408680 547000 1 0 $X=408390 $Y=542790
X673 555 575 561 569 1 5 565 FA1D0BWP7T $T=421560 562680 0 180 $X=408390 $Y=558470
X674 554 549 569 580 1 5 583 FA1D0BWP7T $T=408680 570520 0 0 $X=408390 $Y=570285
X675 227 551 537 542 1 5 566 FA1D0BWP7T $T=421560 586200 1 180 $X=408390 $Y=585965
X676 234 580 566 571 1 5 576 FA1D0BWP7T $T=431080 570520 0 180 $X=417910 $Y=566310
X677 237 588 229 574 1 5 577 FA1D0BWP7T $T=432200 492120 1 180 $X=419030 $Y=491885
X678 558 586 564 592 1 5 241 FA1D0BWP7T $T=419880 507800 1 0 $X=419590 $Y=503590
X679 265 597 577 586 1 5 236 FA1D0BWP7T $T=444520 484280 1 180 $X=431350 $Y=484045
X680 238 246 256 597 1 5 266 FA1D0BWP7T $T=431640 499960 0 0 $X=431350 $Y=499725
X681 18 5 1 15 INVD1BWP7T $T=161720 586200 1 0 $X=161430 $Y=581990
X682 44 5 1 284 INVD1BWP7T $T=186360 515640 0 180 $X=184390 $Y=511430
X683 49 5 1 22 INVD1BWP7T $T=186920 594040 1 180 $X=184950 $Y=593805
X684 50 5 1 33 INVD1BWP7T $T=189720 594040 0 180 $X=187750 $Y=589830
X685 66 5 1 315 INVD1BWP7T $T=208760 523480 0 180 $X=206790 $Y=519270
X686 380 5 1 320 INVD1BWP7T $T=230040 539160 0 180 $X=228070 $Y=534950
X687 85 5 1 332 INVD1BWP7T $T=264760 539160 0 180 $X=262790 $Y=534950
X688 142 5 1 336 INVD1BWP7T $T=313480 554840 0 180 $X=311510 $Y=550630
X689 126 5 1 310 INVD1BWP7T $T=330280 507800 1 180 $X=328310 $Y=507565
X690 182 5 1 168 INVD1BWP7T $T=355480 578360 1 180 $X=353510 $Y=578125
X691 466 5 1 190 INVD1BWP7T $T=367240 515640 0 0 $X=366950 $Y=515405
X692 524 5 1 164 INVD1BWP7T $T=373400 578360 0 180 $X=371430 $Y=574150
X693 232 5 1 181 INVD1BWP7T $T=426600 578360 1 180 $X=424630 $Y=578125
X806 6 5 282 285 1 ND2D1BWP7T $T=156120 492120 0 0 $X=155830 $Y=491885
X807 19 5 293 13 1 ND2D1BWP7T $T=162280 484280 1 180 $X=159750 $Y=484045
X808 6 5 23 16 1 ND2D1BWP7T $T=162280 484280 0 0 $X=161990 $Y=484045
X809 26 5 300 14 1 ND2D1BWP7T $T=167320 507800 0 0 $X=167030 $Y=507565
X810 32 5 303 16 1 ND2D1BWP7T $T=174600 507800 1 180 $X=172070 $Y=507565
X811 36 5 305 319 1 ND2D1BWP7T $T=180200 499960 0 0 $X=179910 $Y=499725
X812 60 5 58 38 1 ND2D1BWP7T $T=205400 531320 0 180 $X=202870 $Y=527110
X813 44 5 384 85 1 ND2D1BWP7T $T=230040 539160 1 0 $X=229750 $Y=534950
X814 426 5 425 379 1 ND2D1BWP7T $T=284920 523480 1 180 $X=282390 $Y=523245
X815 111 5 436 114 1 ND2D1BWP7T $T=282680 531320 1 0 $X=282390 $Y=527110
X816 380 5 429 112 1 ND2D1BWP7T $T=284920 531320 1 180 $X=282390 $Y=531085
X817 119 5 449 426 1 ND2D1BWP7T $T=291640 515640 0 0 $X=291350 $Y=515405
X818 453 5 447 379 1 ND2D1BWP7T $T=300600 562680 1 180 $X=298070 $Y=562445
X819 344 5 419 126 1 ND2D1BWP7T $T=300600 570520 0 180 $X=298070 $Y=566310
X820 66 5 439 142 1 ND2D1BWP7T $T=310680 547000 0 0 $X=310390 $Y=546765
X821 460 5 451 440 1 ND2D1BWP7T $T=318520 515640 1 180 $X=315990 $Y=515405
X822 505 5 511 188 1 ND2D1BWP7T $T=357720 578360 1 0 $X=357430 $Y=574150
X823 524 5 552 219 1 ND2D1BWP7T $T=397480 562680 0 0 $X=397190 $Y=562445
X824 182 5 590 235 1 ND2D1BWP7T $T=429400 594040 0 0 $X=429110 $Y=593805
X825 249 5 593 188 1 ND2D1BWP7T $T=437240 594040 1 180 $X=434710 $Y=593805
X826 250 5 594 505 1 ND2D1BWP7T $T=441160 531320 0 180 $X=438630 $Y=527110
X827 245 5 591 191 1 ND2D1BWP7T $T=442280 554840 1 180 $X=439750 $Y=554605
X828 259 5 599 264 1 ND2D1BWP7T $T=441160 594040 0 0 $X=440870 $Y=593805
X849 46 5 1 335 INVD0BWP7T $T=186920 578360 0 0 $X=186630 $Y=578125
X850 52 5 1 328 INVD0BWP7T $T=188600 586200 1 180 $X=186630 $Y=585965
X851 349 5 1 352 INVD0BWP7T $T=208200 531320 1 180 $X=206230 $Y=531085
X852 358 5 1 356 INVD0BWP7T $T=209880 515640 1 180 $X=207910 $Y=515405
X853 365 5 1 346 INVD0BWP7T $T=217720 539160 1 180 $X=215750 $Y=538925
X854 413 5 1 431 INVD0BWP7T $T=294440 499960 1 180 $X=292470 $Y=499725
X855 427 5 1 406 INVD0BWP7T $T=303400 570520 1 0 $X=303110 $Y=566310
X856 443 5 1 405 INVD0BWP7T $T=314600 499960 1 180 $X=312630 $Y=499725
X857 433 5 1 151 INVD0BWP7T $T=318520 492120 0 180 $X=316550 $Y=487910
X858 474 5 1 467 INVD0BWP7T $T=327480 547000 1 180 $X=325510 $Y=546765
X859 467 5 1 481 INVD0BWP7T $T=335320 547000 1 0 $X=335030 $Y=542790
X860 480 5 1 482 INVD0BWP7T $T=338680 547000 0 180 $X=336710 $Y=542790
X861 154 5 1 490 INVD0BWP7T $T=342040 578360 0 0 $X=341750 $Y=578125
X862 485 5 1 174 INVD0BWP7T $T=347640 499960 1 0 $X=347350 $Y=495750
X863 500 5 1 501 INVD0BWP7T $T=349320 531320 0 0 $X=349030 $Y=531085
X864 502 5 1 503 INVD0BWP7T $T=351000 531320 0 0 $X=350710 $Y=531085
X865 509 5 1 516 INVD0BWP7T $T=358840 539160 0 0 $X=358550 $Y=538925
X866 556 5 1 558 INVD0BWP7T $T=400280 507800 1 0 $X=399990 $Y=503590
X867 361 366 75 364 5 1 OAI21D0BWP7T $T=218280 570520 0 0 $X=217990 $Y=570285
X868 382 418 105 358 5 1 OAI21D0BWP7T $T=269240 507800 0 0 $X=268950 $Y=507565
X869 488 487 160 509 5 1 OAI21D0BWP7T $T=356040 539160 0 0 $X=355750 $Y=538925
X870 507 512 186 171 5 1 OAI21D0BWP7T $T=357720 507800 0 0 $X=357430 $Y=507565
X871 523 522 198 171 5 1 OAI21D0BWP7T $T=384040 507800 1 0 $X=383750 $Y=503590
X872 546 573 557 547 5 1 OAI21D0BWP7T $T=416520 531320 1 180 $X=413430 $Y=531085
X873 572 584 541 171 5 1 OAI21D0BWP7T $T=427720 531320 1 180 $X=424630 $Y=531085
X900 7 5 14 16 1 286 ND3D0BWP7T $T=159480 507800 1 0 $X=159190 $Y=503590
X901 441 5 426 440 1 443 ND3D0BWP7T $T=297240 515640 1 180 $X=294150 $Y=515405
X902 160 5 505 182 1 509 ND3D0BWP7T $T=356040 578360 0 0 $X=355750 $Y=578125
X903 473 5 505 191 1 192 ND3D0BWP7T $T=366680 594040 0 0 $X=366390 $Y=593805
X904 5 1 DCAP16BWP7T $T=156120 507800 0 0 $X=155830 $Y=507565
X905 5 1 DCAP16BWP7T $T=156120 515640 0 0 $X=155830 $Y=515405
X906 5 1 DCAP16BWP7T $T=156120 578360 1 0 $X=155830 $Y=574150
X907 5 1 DCAP16BWP7T $T=166760 570520 0 0 $X=166470 $Y=570285
X908 5 1 DCAP16BWP7T $T=174040 539160 1 0 $X=173750 $Y=534950
X909 5 1 DCAP16BWP7T $T=174040 554840 1 0 $X=173750 $Y=550630
X910 5 1 DCAP16BWP7T $T=174040 562680 1 0 $X=173750 $Y=558470
X911 5 1 DCAP16BWP7T $T=174040 586200 0 0 $X=173750 $Y=585965
X912 5 1 DCAP16BWP7T $T=180760 523480 1 0 $X=180470 $Y=519270
X913 5 1 DCAP16BWP7T $T=180760 570520 0 0 $X=180470 $Y=570285
X914 5 1 DCAP16BWP7T $T=185800 515640 0 0 $X=185510 $Y=515405
X915 5 1 DCAP16BWP7T $T=186920 578360 1 0 $X=186630 $Y=574150
X916 5 1 DCAP16BWP7T $T=188040 554840 1 0 $X=187750 $Y=550630
X917 5 1 DCAP16BWP7T $T=198120 484280 0 0 $X=197830 $Y=484045
X918 5 1 DCAP16BWP7T $T=198120 499960 0 0 $X=197830 $Y=499725
X919 5 1 DCAP16BWP7T $T=211560 492120 1 0 $X=211270 $Y=487910
X920 5 1 DCAP16BWP7T $T=214360 507800 1 0 $X=214070 $Y=503590
X921 5 1 DCAP16BWP7T $T=216040 515640 1 0 $X=215750 $Y=511430
X922 5 1 DCAP16BWP7T $T=216040 539160 1 0 $X=215750 $Y=534950
X923 5 1 DCAP16BWP7T $T=223320 531320 1 0 $X=223030 $Y=527110
X924 5 1 DCAP16BWP7T $T=226680 523480 1 0 $X=226390 $Y=519270
X925 5 1 DCAP16BWP7T $T=227240 562680 1 0 $X=226950 $Y=558470
X926 5 1 DCAP16BWP7T $T=230040 531320 0 0 $X=229750 $Y=531085
X927 5 1 DCAP16BWP7T $T=240120 499960 0 0 $X=239830 $Y=499725
X928 5 1 DCAP16BWP7T $T=240120 515640 0 0 $X=239830 $Y=515405
X929 5 1 DCAP16BWP7T $T=240120 531320 1 0 $X=239830 $Y=527110
X930 5 1 DCAP16BWP7T $T=240120 539160 0 0 $X=239830 $Y=538925
X931 5 1 DCAP16BWP7T $T=240120 554840 0 0 $X=239830 $Y=554605
X932 5 1 DCAP16BWP7T $T=240120 570520 1 0 $X=239830 $Y=566310
X933 5 1 DCAP16BWP7T $T=240120 578360 1 0 $X=239830 $Y=574150
X934 5 1 DCAP16BWP7T $T=258040 507800 0 0 $X=257750 $Y=507565
X935 5 1 DCAP16BWP7T $T=258040 586200 1 0 $X=257750 $Y=581990
X936 5 1 DCAP16BWP7T $T=258600 515640 0 0 $X=258310 $Y=515405
X937 5 1 DCAP16BWP7T $T=263640 594040 1 0 $X=263350 $Y=589830
X938 5 1 DCAP16BWP7T $T=264760 539160 1 0 $X=264470 $Y=534950
X939 5 1 DCAP16BWP7T $T=270920 570520 1 0 $X=270630 $Y=566310
X940 5 1 DCAP16BWP7T $T=271480 515640 0 0 $X=271190 $Y=515405
X941 5 1 DCAP16BWP7T $T=271480 562680 0 0 $X=271190 $Y=562445
X942 5 1 DCAP16BWP7T $T=272040 507800 0 0 $X=271750 $Y=507565
X943 5 1 DCAP16BWP7T $T=282120 499960 0 0 $X=281830 $Y=499725
X944 5 1 DCAP16BWP7T $T=282120 554840 0 0 $X=281830 $Y=554605
X945 5 1 DCAP16BWP7T $T=282120 562680 0 0 $X=281830 $Y=562445
X946 5 1 DCAP16BWP7T $T=282120 570520 1 0 $X=281830 $Y=566310
X947 5 1 DCAP16BWP7T $T=282120 586200 1 0 $X=281830 $Y=581990
X948 5 1 DCAP16BWP7T $T=287720 594040 0 0 $X=287430 $Y=593805
X949 5 1 DCAP16BWP7T $T=300040 547000 0 0 $X=299750 $Y=546765
X950 5 1 DCAP16BWP7T $T=300040 554840 1 0 $X=299750 $Y=550630
X951 5 1 DCAP16BWP7T $T=306760 515640 1 0 $X=306470 $Y=511430
X952 5 1 DCAP16BWP7T $T=310120 523480 0 0 $X=309830 $Y=523245
X953 5 1 DCAP16BWP7T $T=311240 531320 0 0 $X=310950 $Y=531085
X954 5 1 DCAP16BWP7T $T=313480 554840 1 0 $X=313190 $Y=550630
X955 5 1 DCAP16BWP7T $T=313480 562680 1 0 $X=313190 $Y=558470
X956 5 1 DCAP16BWP7T $T=313480 594040 0 0 $X=313190 $Y=593805
X957 5 1 DCAP16BWP7T $T=314040 570520 1 0 $X=313750 $Y=566310
X958 5 1 DCAP16BWP7T $T=324120 499960 1 0 $X=323830 $Y=495750
X959 5 1 DCAP16BWP7T $T=324120 523480 1 0 $X=323830 $Y=519270
X960 5 1 DCAP16BWP7T $T=324120 539160 0 0 $X=323830 $Y=538925
X961 5 1 DCAP16BWP7T $T=331400 531320 1 0 $X=331110 $Y=527110
X962 5 1 DCAP16BWP7T $T=342040 507800 1 0 $X=341750 $Y=503590
X963 5 1 DCAP16BWP7T $T=348200 507800 0 0 $X=347910 $Y=507565
X964 5 1 DCAP16BWP7T $T=348760 515640 0 0 $X=348470 $Y=515405
X965 5 1 DCAP16BWP7T $T=349320 570520 0 0 $X=349030 $Y=570285
X966 5 1 DCAP16BWP7T $T=352120 531320 1 0 $X=351830 $Y=527110
X967 5 1 DCAP16BWP7T $T=352680 586200 1 0 $X=352390 $Y=581990
X968 5 1 DCAP16BWP7T $T=356040 507800 1 0 $X=355750 $Y=503590
X969 5 1 DCAP16BWP7T $T=356040 547000 0 0 $X=355750 $Y=546765
X970 5 1 DCAP16BWP7T $T=366120 499960 0 0 $X=365830 $Y=499725
X971 5 1 DCAP16BWP7T $T=366120 515640 1 0 $X=365830 $Y=511430
X972 5 1 DCAP16BWP7T $T=366120 539160 1 0 $X=365830 $Y=534950
X973 5 1 DCAP16BWP7T $T=372840 578360 0 0 $X=372550 $Y=578125
X974 5 1 DCAP16BWP7T $T=408120 492120 0 0 $X=407830 $Y=491885
X975 5 1 DCAP16BWP7T $T=408120 499960 1 0 $X=407830 $Y=495750
X976 5 1 DCAP16BWP7T $T=408120 507800 1 0 $X=407830 $Y=503590
X977 5 1 DCAP16BWP7T $T=408120 523480 1 0 $X=407830 $Y=519270
X978 5 1 DCAP16BWP7T $T=408120 554840 1 0 $X=407830 $Y=550630
X979 5 1 DCAP16BWP7T $T=408120 570520 1 0 $X=407830 $Y=566310
X980 5 1 DCAP16BWP7T $T=421560 484280 0 0 $X=421270 $Y=484045
X981 5 1 DCAP16BWP7T $T=421560 499960 0 0 $X=421270 $Y=499725
X982 5 1 DCAP16BWP7T $T=426040 547000 0 0 $X=425750 $Y=546765
X983 5 1 DCAP16BWP7T $T=431080 523480 1 0 $X=430790 $Y=519270
X984 5 1 DCAP16BWP7T $T=432760 507800 1 0 $X=432470 $Y=503590
X985 5 1 DCAP16BWP7T $T=437800 492120 0 0 $X=437510 $Y=491885
X986 5 1 DCAP16BWP7T $T=439480 562680 1 0 $X=439190 $Y=558470
X987 5 1 DCAP16BWP7T $T=439480 570520 0 0 $X=439190 $Y=570285
X1033 316 5 326 406 396 1 NR3D1BWP7T $T=258600 515640 1 180 $X=253830 $Y=515405
X1034 173 5 166 490 495 1 NR3D1BWP7T $T=351000 570520 1 0 $X=350710 $Y=566310
X1035 61 346 5 1 347 349 MAOI222D1BWP7T $T=206520 531320 1 180 $X=201750 $Y=531085
X1036 143 140 5 1 141 138 MAOI222D1BWP7T $T=313480 594040 1 180 $X=308710 $Y=593805
X1037 159 468 5 1 477 474 MAOI222D1BWP7T $T=335880 570520 0 180 $X=331110 $Y=566310
X1038 501 508 5 1 478 502 MAOI222D1BWP7T $T=356040 531320 0 0 $X=355750 $Y=531085
X1039 541 562 5 1 568 556 MAOI222D1BWP7T $T=415400 515640 0 180 $X=410630 $Y=511430
X1040 48 47 5 324 333 1 AOI21D1BWP7T $T=189720 586200 0 180 $X=186070 $Y=581990
X1041 406 425 5 396 409 1 AOI21D1BWP7T $T=269240 515640 1 0 $X=268950 $Y=511430
X1042 490 511 5 495 477 1 AOI21D1BWP7T $T=366680 562680 0 0 $X=366390 $Y=562445
X1043 490 511 5 495 471 1 AOI21D1BWP7T $T=368360 570520 1 0 $X=368070 $Y=566310
X1044 198 523 5 522 197 1 AOI21D1BWP7T $T=375080 499960 0 180 $X=371430 $Y=495750
X1045 285 11 1 5 INVD2BWP7T $T=157800 484280 0 0 $X=157510 $Y=484045
X1046 426 326 1 5 INVD2BWP7T $T=271480 515640 1 180 $X=268950 $Y=515405
X1047 111 318 1 5 INVD2BWP7T $T=285480 492120 0 180 $X=282950 $Y=487910
X1048 440 42 1 5 INVD2BWP7T $T=286040 523480 0 180 $X=283510 $Y=519270
X1049 145 127 1 5 INVD2BWP7T $T=315160 547000 1 180 $X=312630 $Y=546765
X1050 505 166 1 5 INVD2BWP7T $T=358280 570520 1 0 $X=357990 $Y=566310
X1051 188 173 1 5 INVD2BWP7T $T=382360 578360 1 0 $X=382070 $Y=574150
X1052 218 176 1 5 INVD2BWP7T $T=399720 562680 0 180 $X=397190 $Y=558470
X1099 9 302 5 1 294 DFQD0BWP7T $T=169560 554840 0 0 $X=169270 $Y=554605
X1100 9 308 5 1 342 DFQD0BWP7T $T=181880 554840 0 0 $X=181590 $Y=554605
X1101 9 309 5 1 18 DFQD0BWP7T $T=209320 562680 0 180 $X=198390 $Y=558470
X1102 83 350 5 1 77 DFQD0BWP7T $T=232840 594040 1 180 $X=221910 $Y=593805
X1103 83 392 5 1 89 DFQD0BWP7T $T=251320 594040 0 180 $X=240390 $Y=589830
X1104 83 442 5 1 416 DFQD0BWP7T $T=293320 578360 0 180 $X=282390 $Y=574150
X1105 83 444 5 1 427 DFQD0BWP7T $T=293880 586200 1 180 $X=282950 $Y=585965
X1106 9 458 5 1 441 DFQD0BWP7T $T=308440 515640 1 180 $X=297510 $Y=515405
X1107 9 450 5 1 452 DFQD0BWP7T $T=309560 539160 1 180 $X=298630 $Y=538925
X1108 9 139 5 1 454 DFQD0BWP7T $T=312920 492120 0 180 $X=301990 $Y=487910
X1109 9 149 5 1 459 DFQD0BWP7T $T=318520 507800 0 180 $X=307590 $Y=503590
X1110 9 146 5 1 460 DFQD0BWP7T $T=318520 523480 0 180 $X=307590 $Y=519270
X1111 83 465 5 1 461 DFQD0BWP7T $T=318520 594040 0 180 $X=307590 $Y=589830
X1112 9 475 5 1 153 DFQD0BWP7T $T=335320 515640 1 180 $X=324390 $Y=515405
X1113 9 469 5 1 160 DFQD0BWP7T $T=324680 547000 1 0 $X=324390 $Y=542790
X1114 83 470 5 1 473 DFQD0BWP7T $T=324680 570520 0 0 $X=324390 $Y=570285
X1115 83 463 5 1 154 DFQD0BWP7T $T=335320 586200 0 180 $X=324390 $Y=581990
X1116 9 476 5 1 155 DFQD0BWP7T $T=336440 499960 1 180 $X=325510 $Y=499725
X1117 9 492 5 1 163 DFQD0BWP7T $T=347640 523480 0 180 $X=336710 $Y=519270
X1118 9 493 5 1 466 DFQD0BWP7T $T=348200 507800 1 180 $X=337270 $Y=507565
X1119 9 504 5 1 485 DFQD0BWP7T $T=359960 492120 1 180 $X=349030 $Y=491885
X1120 9 529 5 1 207 DFQD0BWP7T $T=375640 515640 1 0 $X=375350 $Y=511430
X1121 9 550 5 1 201 DFQD0BWP7T $T=391880 523480 0 0 $X=391590 $Y=523245
X1122 222 570 5 1 218 DFQD0BWP7T $T=408680 531320 1 0 $X=408390 $Y=527110
X1123 222 581 5 1 226 DFQD0BWP7T $T=431080 523480 0 180 $X=420150 $Y=519270
X1124 222 253 5 1 235 DFQD0BWP7T $T=443400 531320 1 180 $X=432470 $Y=531085
X1125 171 144 5 1 INVD4BWP7T $T=344280 586200 1 180 $X=340070 $Y=585965
X1126 48 5 1 45 25 324 NR3D0BWP7T $T=188040 594040 0 180 $X=184950 $Y=589830
X1127 507 493 186 512 5 1 AOI21D0BWP7T $T=357720 515640 1 0 $X=357430 $Y=511430
X1128 572 581 541 584 5 1 AOI21D0BWP7T $T=419880 531320 0 0 $X=419590 $Y=531085
X1129 14 16 5 1 283 AN2D1BWP7T $T=162840 507800 1 0 $X=162550 $Y=503590
X1130 14 31 5 1 29 AN2D1BWP7T $T=172360 507800 1 180 $X=169270 $Y=507565
X1131 32 31 5 1 304 AN2D1BWP7T $T=171240 484280 0 0 $X=170950 $Y=484045
X1132 34 36 5 1 306 AN2D1BWP7T $T=174040 484280 0 0 $X=173750 $Y=484045
X1133 34 38 5 1 39 AN2D1BWP7T $T=177400 499960 0 0 $X=177110 $Y=499725
X1134 319 38 5 1 348 AN2D1BWP7T $T=200920 523480 1 0 $X=200630 $Y=519270
X1135 114 426 5 1 422 AN2D1BWP7T $T=287720 531320 1 180 $X=284630 $Y=531085
X1136 133 130 5 1 430 AN2D1BWP7T $T=301720 586200 1 180 $X=298630 $Y=585965
X1137 453 131 5 1 128 AN2D1BWP7T $T=302280 547000 0 180 $X=299190 $Y=542790
X1138 453 440 5 1 428 AN2D1BWP7T $T=311240 531320 1 180 $X=308150 $Y=531085
X1139 460 131 5 1 137 AN2D1BWP7T $T=311240 578360 0 180 $X=308150 $Y=574150
X1140 180 131 5 1 464 AN2D1BWP7T $T=351560 578360 1 180 $X=348470 $Y=578125
X1141 540 171 5 1 529 AN2D1BWP7T $T=389640 507800 0 180 $X=386550 $Y=503590
X1142 220 505 5 1 561 AN2D1BWP7T $T=399720 562680 1 0 $X=399430 $Y=558470
X1143 245 131 5 1 240 AN2D1BWP7T $T=434440 594040 1 180 $X=431350 $Y=593805
X1144 249 191 5 1 575 AN2D1BWP7T $T=440040 554840 1 180 $X=436950 $Y=554605
X1145 592 171 5 1 598 AN2D1BWP7T $T=441720 523480 1 0 $X=441430 $Y=519270
X1146 347 61 365 1 5 369 XOR3D0BWP7T $T=212120 547000 1 0 $X=211830 $Y=542790
X1147 87 101 433 1 5 109 XOR3D0BWP7T $T=267000 484280 0 0 $X=266710 $Y=484045
X1148 508 478 500 1 5 518 XOR3D0BWP7T $T=377880 507800 0 180 $X=368070 $Y=503590
X1149 361 364 75 1 5 367 XNR3D0BWP7T $T=211560 586200 1 0 $X=211270 $Y=581990
X1150 405 409 417 1 5 420 XNR3D0BWP7T $T=255800 515640 1 0 $X=255510 $Y=511430
X1151 97 81 82 1 5 421 XNR3D0BWP7T $T=255800 578360 0 0 $X=255510 $Y=578125
X1152 96 103 93 1 5 124 XNR3D0BWP7T $T=288280 492120 1 0 $X=287990 $Y=487910
X1153 159 471 468 1 5 462 XNR3D0BWP7T $T=334200 554840 1 180 $X=324390 $Y=554605
X1154 546 547 557 1 5 560 XNR3D0BWP7T $T=393000 539160 1 0 $X=392710 $Y=534950
X1155 361 75 5 390 366 1 IOA21D0BWP7T $T=266440 570520 0 0 $X=266150 $Y=570285
X1156 71 150 5 458 448 1 IOA21D0BWP7T $T=318520 492120 1 180 $X=314870 $Y=491885
X1157 152 473 5 158 157 1 IOA21D0BWP7T $T=333080 586200 1 180 $X=329430 $Y=585965
X1158 152 485 5 470 486 1 IOA21D0BWP7T $T=338120 578360 1 0 $X=337830 $Y=574150
X1159 546 557 5 567 573 1 IOA21D0BWP7T $T=420440 554840 1 0 $X=420150 $Y=550630
X1160 258 261 5 263 269 1 IOA21D0BWP7T $T=441160 586200 0 0 $X=440870 $Y=585965
X1161 443 5 65 441 1 438 448 OAI211D0BWP7T $T=289960 515640 1 0 $X=289670 $Y=511430
X1162 192 5 171 473 1 517 486 OAI211D0BWP7T $T=370040 586200 1 180 $X=366390 $Y=585965
X1163 59 65 355 71 5 1 350 AO22D0BWP7T $T=209880 578360 0 180 $X=205110 $Y=574150
X1164 86 65 381 71 5 1 80 AO22D0BWP7T $T=232840 578360 0 180 $X=228070 $Y=574150
X1165 125 65 432 71 5 1 450 AO22D0BWP7T $T=298920 507800 0 180 $X=294150 $Y=503590
X1166 207 171 544 152 5 1 536 AO22D0BWP7T $T=400280 507800 0 180 $X=395510 $Y=503590
X1167 243 171 579 152 5 1 248 AO22D0BWP7T $T=441160 515640 0 180 $X=436390 $Y=511430
X1168 97 82 81 375 5 1 MAOI222D2BWP7T $T=233400 586200 1 180 $X=225830 $Y=585965
X1169 405 417 409 423 5 1 MAOI222D2BWP7T $T=289960 507800 0 180 $X=282390 $Y=503590
X1170 9 288 5 1 13 DFQD1BWP7T $T=156120 523480 1 0 $X=155830 $Y=519270
X1171 9 287 5 1 24 DFQD1BWP7T $T=156120 570520 0 0 $X=155830 $Y=570285
X1172 9 281 5 1 27 DFQD1BWP7T $T=156680 554840 0 0 $X=156390 $Y=554605
X1173 9 289 5 1 285 DFQD1BWP7T $T=157240 531320 0 0 $X=156950 $Y=531085
X1174 9 290 5 1 31 DFQD1BWP7T $T=167320 547000 1 0 $X=167030 $Y=542790
X1175 9 298 5 1 26 DFQD1BWP7T $T=167880 523480 1 0 $X=167590 $Y=519270
X1176 9 301 5 1 34 DFQD1BWP7T $T=170120 531320 0 0 $X=169830 $Y=531085
X1177 9 337 5 1 49 DFQD1BWP7T $T=203160 570520 1 0 $X=202870 $Y=566310
X1178 9 91 5 1 327 DFQD1BWP7T $T=251320 484280 1 180 $X=240390 $Y=484045
X1179 83 411 5 1 95 DFQD1BWP7T $T=263640 594040 0 180 $X=252710 $Y=589830
X1180 83 430 5 1 319 DFQD1BWP7T $T=276520 594040 1 180 $X=265590 $Y=593805
X1181 83 456 5 1 379 DFQD1BWP7T $T=306760 578360 0 180 $X=295830 $Y=574150
X1182 9 457 5 1 426 DFQD1BWP7T $T=308440 499960 1 180 $X=297510 $Y=499725
X1183 9 147 5 1 453 DFQD1BWP7T $T=318520 539160 0 180 $X=307590 $Y=534950
X1184 83 464 5 1 119 DFQD1BWP7T $T=318520 562680 1 180 $X=307590 $Y=562445
X1185 83 148 5 1 114 DFQD1BWP7T $T=318520 578360 1 180 $X=307590 $Y=578125
X1186 9 491 5 1 479 DFQD1BWP7T $T=347640 499960 0 180 $X=336710 $Y=495750
X1187 9 506 5 1 175 DFQD1BWP7T $T=360520 523480 0 180 $X=349590 $Y=519270
X1188 9 519 5 1 505 DFQD1BWP7T $T=366680 523480 0 0 $X=366390 $Y=523245
X1189 9 536 5 1 196 DFQD1BWP7T $T=387960 523480 1 180 $X=377030 $Y=523245
X1190 9 545 5 1 524 DFQD1BWP7T $T=389080 515640 1 0 $X=388790 $Y=511430
X1191 222 598 5 1 243 DFQD1BWP7T $T=443400 515640 1 180 $X=432470 $Y=515405
X1192 71 84 5 1 369 392 79 MOAI22D0BWP7T $T=258040 578360 0 180 $X=253830 $Y=574150
X1193 71 427 5 1 79 104 421 MOAI22D0BWP7T $T=272600 578360 1 180 $X=268390 $Y=578125
X1194 71 105 5 1 398 411 79 MOAI22D0BWP7T $T=273720 570520 1 180 $X=269510 $Y=570285
X1195 71 441 5 1 79 113 110 MOAI22D0BWP7T $T=286600 570520 1 180 $X=282390 $Y=570285
X1196 152 466 5 1 144 463 462 MOAI22D0BWP7T $T=317400 554840 1 180 $X=313190 $Y=554605
X1197 152 177 5 1 499 469 144 MOAI22D0BWP7T $T=352120 531320 0 180 $X=347910 $Y=527110
X1198 152 200 5 1 518 506 144 MOAI22D0BWP7T $T=378440 531320 0 180 $X=374230 $Y=527110
X1199 286 303 67 299 340 5 1 XNR4D0BWP7T $T=201480 507800 1 0 $X=201190 $Y=503590
X1200 437 439 445 446 407 5 1 XNR4D0BWP7T $T=282680 547000 1 0 $X=282390 $Y=542790
X1201 120 447 437 424 415 5 1 XNR4D0BWP7T $T=295560 562680 0 180 $X=282390 $Y=558470
X1202 595 242 589 587 585 5 1 XNR4D0BWP7T $T=436120 554840 1 180 $X=422950 $Y=554605
X1203 233 593 595 596 255 5 1 XNR4D0BWP7T $T=428840 586200 1 0 $X=428550 $Y=581990
X1204 115 8 5 1 BUFFD12BWP7T $T=343160 531320 1 180 $X=330550 $Y=531085
X1205 305 300 299 293 282 5 1 XOR4D0BWP7T $T=175720 499960 0 180 $X=162550 $Y=495750
X1206 357 70 72 73 76 5 1 XOR4D0BWP7T $T=208200 484280 0 0 $X=207910 $Y=484045
X1207 399 402 407 410 416 5 1 XOR4D0BWP7T $T=251320 570520 1 0 $X=251030 $Y=566310
X1208 436 429 424 384 419 5 1 XOR4D0BWP7T $T=276520 539160 1 180 $X=263350 $Y=538925
X1209 449 451 446 435 414 5 1 XOR4D0BWP7T $T=301160 531320 0 180 $X=287990 $Y=527110
X1210 565 559 585 576 231 5 1 XOR4D0BWP7T $T=414280 586200 1 0 $X=413990 $Y=581990
X1211 594 591 587 582 583 5 1 XOR4D0BWP7T $T=434440 547000 0 180 $X=421270 $Y=542790
X1212 239 590 596 552 599 5 1 XOR4D0BWP7T $T=431080 570520 1 0 $X=430790 $Y=566310
X1213 344 5 1 307 CKND1BWP7T $T=191960 570520 0 180 $X=189990 $Y=566310
X1214 201 5 1 538 CKND1BWP7T $T=386840 578360 1 0 $X=386550 $Y=574150
X1215 30 28 5 1 BUFFD1P5BWP7T $T=170680 578360 0 180 $X=167590 $Y=574150
X1216 479 161 5 1 BUFFD1P5BWP7T $T=334200 499960 1 0 $X=333910 $Y=495750
X1217 204 205 1 206 5 208 523 AOI22D1BWP7T $T=382920 499960 0 0 $X=382630 $Y=499725
X1218 294 5 1 21 CKBD1BWP7T $T=160600 594040 1 0 $X=160310 $Y=589830
X1219 342 5 1 56 CKBD1BWP7T $T=190280 562680 1 0 $X=189990 $Y=558470
X1220 122 5 1 380 CKBD1BWP7T $T=296120 570520 0 180 $X=293590 $Y=566310
X1221 452 5 1 86 CKBD1BWP7T $T=296680 539160 0 0 $X=296390 $Y=538925
X1222 459 5 1 112 CKBD1BWP7T $T=305640 507800 1 0 $X=305350 $Y=503590
X1223 461 5 1 440 CKBD1BWP7T $T=314040 570520 0 180 $X=311510 $Y=566310
X1224 454 5 1 344 CKBD1BWP7T $T=333640 492120 1 180 $X=331110 $Y=491885
X1225 538 5 1 172 CKBD1BWP7T $T=384600 578360 1 0 $X=384310 $Y=574150
X1226 252 5 1 250 CKBD1BWP7T $T=440600 547000 1 180 $X=438070 $Y=546765
X1227 379 316 5 1 INVD1P5BWP7T $T=270920 570520 0 180 $X=268390 $Y=566310
X1228 189 187 1 5 187 507 189 MAOI22D0BWP7T $T=367240 492120 0 0 $X=366950 $Y=491885
X1229 562 568 1 5 568 572 562 MAOI22D0BWP7T $T=408680 515640 0 0 $X=408390 $Y=515405
X1230 7 283 286 1 5 295 OA21D0BWP7T $T=156120 499960 1 0 $X=155830 $Y=495750
X1231 5 1 ICV_76 $T=155000 492120 1 0 $X=154710 $Y=487910
X1232 5 1 ICV_76 $T=155000 499960 0 0 $X=154710 $Y=499725
X1233 5 1 ICV_76 $T=155000 531320 1 0 $X=154710 $Y=527110
X1234 5 1 ICV_76 $T=155000 539160 1 0 $X=154710 $Y=534950
X1235 5 1 ICV_76 $T=155000 539160 0 0 $X=154710 $Y=538925
X1236 5 1 ICV_76 $T=155000 554840 1 0 $X=154710 $Y=550630
X1237 5 1 ICV_76 $T=155000 562680 1 0 $X=154710 $Y=558470
X1238 5 1 ICV_76 $T=155000 586200 0 0 $X=154710 $Y=585965
X1239 5 1 ICV_76 $T=197000 539160 1 0 $X=196710 $Y=534950
X1240 5 1 ICV_76 $T=197000 539160 0 0 $X=196710 $Y=538925
X1241 5 1 ICV_76 $T=197000 562680 0 0 $X=196710 $Y=562445
X1242 5 1 ICV_76 $T=197000 594040 0 0 $X=196710 $Y=593805
X1243 5 1 ICV_76 $T=239000 570520 0 0 $X=238710 $Y=570285
X1244 5 1 ICV_76 $T=239000 586200 1 0 $X=238710 $Y=581990
X1245 5 1 ICV_76 $T=239000 594040 0 0 $X=238710 $Y=593805
X1246 5 1 ICV_76 $T=281000 554840 1 0 $X=280710 $Y=550630
X1247 5 1 ICV_76 $T=281000 578360 0 0 $X=280710 $Y=578125
X1248 5 1 ICV_76 $T=281000 594040 1 0 $X=280710 $Y=589830
X1249 5 1 ICV_76 $T=365000 547000 0 0 $X=364710 $Y=546765
X1250 5 1 ICV_76 $T=407000 594040 0 0 $X=406710 $Y=593805
X1251 5 1 ICV_41 $T=163960 578360 0 0 $X=163670 $Y=578125
X1252 5 1 ICV_41 $T=198120 586200 1 0 $X=197830 $Y=581990
X1253 5 1 ICV_41 $T=211560 586200 0 0 $X=211270 $Y=585965
X1254 5 1 ICV_41 $T=266440 554840 1 0 $X=266150 $Y=550630
X1255 5 1 ICV_41 $T=282120 539160 0 0 $X=281830 $Y=538925
X1256 5 1 ICV_41 $T=309000 499960 1 0 $X=308710 $Y=495750
X1257 5 1 ICV_41 $T=309560 539160 0 0 $X=309270 $Y=538925
X1258 5 1 ICV_41 $T=333640 492120 0 0 $X=333350 $Y=491885
X1259 5 1 ICV_41 $T=349880 562680 0 0 $X=349590 $Y=562445
X1260 5 1 ICV_41 $T=384040 562680 1 0 $X=383750 $Y=558470
X1261 5 1 ICV_41 $T=392440 554840 1 0 $X=392150 $Y=550630
X1262 5 1 ICV_41 $T=393000 492120 1 0 $X=392710 $Y=487910
X1263 5 1 ICV_41 $T=393000 499960 1 0 $X=392710 $Y=495750
X1264 5 1 ICV_41 $T=393560 570520 1 0 $X=393270 $Y=566310
X1265 5 1 ICV_41 $T=408120 554840 0 0 $X=407830 $Y=554605
X1266 5 1 ICV_41 $T=408120 578360 0 0 $X=407830 $Y=578125
X1267 5 1 ICV_41 $T=426040 578360 1 0 $X=425750 $Y=574150
X1268 5 1 ICV_37 $T=156120 507800 1 0 $X=155830 $Y=503590
X1269 5 1 ICV_37 $T=156120 586200 1 0 $X=155830 $Y=581990
X1270 5 1 ICV_37 $T=156120 594040 0 0 $X=155830 $Y=593805
X1271 5 1 ICV_37 $T=166760 562680 0 0 $X=166470 $Y=562445
X1272 5 1 ICV_37 $T=174040 499960 0 0 $X=173750 $Y=499725
X1273 5 1 ICV_37 $T=181880 594040 0 0 $X=181590 $Y=593805
X1274 5 1 ICV_37 $T=183000 539160 1 0 $X=182710 $Y=534950
X1275 5 1 ICV_37 $T=193640 499960 1 0 $X=193350 $Y=495750
X1276 5 1 ICV_37 $T=198120 507800 1 0 $X=197830 $Y=503590
X1277 5 1 ICV_37 $T=227800 499960 0 0 $X=227510 $Y=499725
X1278 5 1 ICV_37 $T=235640 523480 1 0 $X=235350 $Y=519270
X1279 5 1 ICV_37 $T=235640 539160 0 0 $X=235350 $Y=538925
X1280 5 1 ICV_37 $T=282120 594040 0 0 $X=281830 $Y=593805
X1281 5 1 ICV_37 $T=294440 499960 0 0 $X=294150 $Y=499725
X1282 5 1 ICV_37 $T=303960 523480 1 0 $X=303670 $Y=519270
X1283 5 1 ICV_37 $T=312920 492120 1 0 $X=312630 $Y=487910
X1284 5 1 ICV_37 $T=319640 547000 0 0 $X=319350 $Y=546765
X1285 5 1 ICV_37 $T=319640 586200 0 0 $X=319350 $Y=585965
X1286 5 1 ICV_37 $T=361640 586200 1 0 $X=361350 $Y=581990
X1287 5 1 ICV_37 $T=373400 492120 0 0 $X=373110 $Y=491885
X1288 5 1 ICV_37 $T=394120 562680 0 0 $X=393830 $Y=562445
X1289 5 1 ICV_37 $T=403640 578360 0 0 $X=403350 $Y=578125
X1290 5 1 ICV_37 $T=417080 523480 1 0 $X=416790 $Y=519270
X1291 5 1 ICV_37 $T=417080 554840 1 0 $X=416790 $Y=550630
X1292 5 1 ICV_37 $T=434440 547000 1 0 $X=434150 $Y=542790
X1293 5 1 ICV_37 $T=435000 547000 0 0 $X=434710 $Y=546765
X1294 5 1 ICV_60 $T=174040 539160 0 0 $X=173750 $Y=538925
X1295 5 1 ICV_60 $T=181320 586200 1 0 $X=181030 $Y=581990
X1296 5 1 ICV_60 $T=198120 531320 1 0 $X=197830 $Y=527110
X1297 5 1 ICV_60 $T=198120 570520 1 0 $X=197830 $Y=566310
X1298 5 1 ICV_60 $T=205400 531320 1 0 $X=205110 $Y=527110
X1299 5 1 ICV_60 $T=225000 515640 1 0 $X=224710 $Y=511430
X1300 5 1 ICV_60 $T=249080 515640 0 0 $X=248790 $Y=515405
X1301 5 1 ICV_60 $T=249080 578360 1 0 $X=248790 $Y=574150
X1302 5 1 ICV_60 $T=293880 586200 0 0 $X=293590 $Y=585965
X1303 5 1 ICV_60 $T=324120 492120 1 0 $X=323830 $Y=487910
X1304 5 1 ICV_60 $T=375080 539160 1 0 $X=374790 $Y=534950
X1305 5 1 ICV_60 $T=443960 492120 1 0 $X=443670 $Y=487910
X1306 5 1 ICV_60 $T=443960 507800 0 0 $X=443670 $Y=507565
X1307 5 1 ICV_60 $T=443960 523480 0 0 $X=443670 $Y=523245
X1308 5 1 ICV_60 $T=443960 539160 1 0 $X=443670 $Y=534950
X1309 5 1 ICV_60 $T=443960 539160 0 0 $X=443670 $Y=538925
X1310 5 1 ICV_60 $T=443960 562680 0 0 $X=443670 $Y=562445
X1311 5 1 ICV_60 $T=443960 570520 1 0 $X=443670 $Y=566310
X1312 5 1 ICV_60 $T=443960 594040 1 0 $X=443670 $Y=589830
X1313 5 1 ICV_43 $T=156120 547000 1 0 $X=155830 $Y=542790
X1314 5 1 ICV_43 $T=165080 578360 1 0 $X=164790 $Y=574150
X1315 5 1 ICV_43 $T=176280 515640 1 0 $X=175990 $Y=511430
X1316 5 1 ICV_43 $T=183000 554840 1 0 $X=182710 $Y=550630
X1317 5 1 ICV_43 $T=198120 523480 1 0 $X=197830 $Y=519270
X1318 5 1 ICV_43 $T=226120 515640 0 0 $X=225830 $Y=515405
X1319 5 1 ICV_43 $T=267000 586200 1 0 $X=266710 $Y=581990
X1320 5 1 ICV_43 $T=285480 492120 1 0 $X=285190 $Y=487910
X1321 5 1 ICV_43 $T=291080 570520 1 0 $X=290790 $Y=566310
X1322 5 1 ICV_43 $T=300600 570520 1 0 $X=300310 $Y=566310
X1323 5 1 ICV_43 $T=302840 523480 0 0 $X=302550 $Y=523245
X1324 5 1 ICV_43 $T=305080 562680 0 0 $X=304790 $Y=562445
X1325 5 1 ICV_43 $T=305640 531320 0 0 $X=305350 $Y=531085
X1326 5 1 ICV_43 $T=309000 554840 1 0 $X=308710 $Y=550630
X1327 5 1 ICV_43 $T=366120 578360 1 0 $X=365830 $Y=574150
X1328 5 1 ICV_43 $T=408120 515640 1 0 $X=407830 $Y=511430
X1329 5 1 ICV_43 $T=417080 507800 1 0 $X=416790 $Y=503590
X1330 320 1 8 54 5 NR2XD0BWP7T $T=191960 523480 0 180 $X=189430 $Y=519270
X1331 5 1 ICV_38 $T=192520 507800 0 0 $X=192230 $Y=507565
X1332 5 1 ICV_38 $T=192520 515640 1 0 $X=192230 $Y=511430
X1333 5 1 ICV_38 $T=192520 531320 1 0 $X=192230 $Y=527110
X1334 5 1 ICV_38 $T=192520 570520 0 0 $X=192230 $Y=570285
X1335 5 1 ICV_38 $T=234520 492120 1 0 $X=234230 $Y=487910
X1336 5 1 ICV_38 $T=276520 515640 1 0 $X=276230 $Y=511430
X1337 5 1 ICV_38 $T=276520 539160 0 0 $X=276230 $Y=538925
X1338 5 1 ICV_38 $T=276520 554840 0 0 $X=276230 $Y=554605
X1339 5 1 ICV_38 $T=276520 594040 0 0 $X=276230 $Y=593805
X1340 5 1 ICV_38 $T=318520 492120 1 0 $X=318230 $Y=487910
X1341 5 1 ICV_38 $T=318520 492120 0 0 $X=318230 $Y=491885
X1342 5 1 ICV_38 $T=318520 507800 1 0 $X=318230 $Y=503590
X1343 5 1 ICV_38 $T=318520 523480 1 0 $X=318230 $Y=519270
X1344 5 1 ICV_38 $T=318520 539160 1 0 $X=318230 $Y=534950
X1345 5 1 ICV_38 $T=318520 562680 0 0 $X=318230 $Y=562445
X1346 5 1 ICV_38 $T=318520 578360 0 0 $X=318230 $Y=578125
X1347 5 1 ICV_38 $T=318520 594040 1 0 $X=318230 $Y=589830
X1348 5 1 ICV_38 $T=360520 499960 0 0 $X=360230 $Y=499725
X1349 5 1 ICV_38 $T=360520 515640 1 0 $X=360230 $Y=511430
X1350 5 1 ICV_38 $T=360520 523480 1 0 $X=360230 $Y=519270
X1351 5 1 ICV_38 $T=360520 531320 0 0 $X=360230 $Y=531085
X1352 5 1 ICV_38 $T=360520 539160 0 0 $X=360230 $Y=538925
X1353 5 1 ICV_38 $T=360520 547000 1 0 $X=360230 $Y=542790
X1354 5 1 ICV_38 $T=360520 554840 0 0 $X=360230 $Y=554605
X1355 5 1 ICV_38 $T=360520 570520 1 0 $X=360230 $Y=566310
X1356 5 1 ICV_38 $T=402520 492120 0 0 $X=402230 $Y=491885
X1357 5 1 ICV_38 $T=402520 547000 0 0 $X=402230 $Y=546765
X1358 59 323 5 1 353 354 IAO21D0BWP7T $T=204840 515640 0 0 $X=204550 $Y=515405
X1359 84 383 5 1 362 378 IAO21D0BWP7T $T=232280 515640 1 180 $X=228630 $Y=515405
X1360 175 498 5 1 513 514 IAO21D0BWP7T $T=357160 547000 1 0 $X=356870 $Y=542790
X1361 196 526 5 1 527 521 IAO21D0BWP7T $T=373400 562680 0 0 $X=373110 $Y=562445
X1362 226 247 5 1 238 588 IAO21D0BWP7T $T=437800 492120 1 180 $X=434150 $Y=491885
X1363 379 44 59 1 5 353 AN3D1BWP7T $T=229480 523480 1 180 $X=225830 $Y=523245
X1364 379 66 84 1 5 362 AN3D1BWP7T $T=233960 507800 0 180 $X=230310 $Y=503590
X1365 379 344 327 1 5 334 AN3D1BWP7T $T=266440 554840 0 180 $X=262790 $Y=550630
X1366 188 524 196 1 5 527 AN3D1BWP7T $T=380120 562680 1 180 $X=376470 $Y=562445
X1367 188 201 175 1 5 513 AN3D1BWP7T $T=380120 578360 0 180 $X=376470 $Y=574150
X1368 9 297 16 5 1 DFQD2BWP7T $T=192520 531320 0 180 $X=181030 $Y=527110
X1369 184 1 115 5 171 NR2XD3BWP7T $T=357720 594040 0 180 $X=349030 $Y=589830
X1370 71 327 5 79 78 367 1 MOAI22D1BWP7T $T=228360 578360 0 180 $X=223590 $Y=574150
X1371 71 135 5 79 444 420 1 MOAI22D1BWP7T $T=303960 492120 0 0 $X=303670 $Y=491885
X1372 71 136 5 79 442 445 1 MOAI22D1BWP7T $T=310120 523480 1 180 $X=305350 $Y=523245
X1373 152 226 5 144 225 560 1 MOAI22D1BWP7T $T=424360 515640 1 180 $X=419590 $Y=515405
X1374 152 251 5 144 257 589 1 MOAI22D1BWP7T $T=437800 547000 1 0 $X=437510 $Y=542790
X1375 144 1 187 185 5 504 174 AOI211D1BWP7T $T=360520 499960 1 180 $X=356870 $Y=499725
X1376 8 51 332 1 5 NR2D1P5BWP7T $T=191960 499960 1 180 $X=187750 $Y=499725
X1377 327 314 1 334 339 5 IAO21D1BWP7T $T=186360 539160 0 0 $X=186070 $Y=538925
X1378 71 416 107 106 1 79 5 IOA22D2BWP7T $T=275960 586200 0 180 $X=269510 $Y=581990
X1379 118 9 5 1 INVD10BWP7T $T=291080 499960 0 180 $X=282390 $Y=495750
X1380 8 71 121 5 1 INR2XD4BWP7T $T=307880 554840 1 180 $X=294710 $Y=554605
X1381 86 5 112 379 1 120 ND3D1BWP7T $T=298360 586200 0 180 $X=294710 $Y=581990
X1382 105 5 426 380 1 358 ND3D1BWP7T $T=299480 547000 0 180 $X=295830 $Y=542790
.ENDS
***************************************
.SUBCKT ICV_75 1 2
** N=2 EP=2 IP=4 FDC=12
*.SEEDPROM
X0 2 1 DCAPBWP7T $T=6720 0 0 0 $X=6430 $Y=-235
X1 1 2 ICV_40 $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_74 1 2
** N=2 EP=2 IP=4 FDC=8
*.SEEDPROM
X0 2 1 DCAPBWP7T $T=4480 0 0 0 $X=4190 $Y=-235
X1 1 2 DCAP8BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT OAI21D1BWP7T A1 A2 VDD B ZN VSS
** N=8 EP=6 IP=0 FDC=6
*.SEEDPROM
M0 ZN A1 7 VSS N L=1.8e-07 W=1e-06 $X=760 $Y=345 $D=0
M1 7 A2 ZN VSS N L=1.8e-07 W=1e-06 $X=1480 $Y=345 $D=0
M2 VSS B 7 VSS N L=1.8e-07 W=1e-06 $X=2200 $Y=345 $D=0
M3 8 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=760 $Y=2205 $D=16
M4 VDD A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=1480 $Y=2205 $D=16
M5 ZN B VDD VDD P L=1.8e-07 W=1.37e-06 $X=2200 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_50
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_77
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_78 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215
** N=678 EP=214 IP=4890 FDC=13216
*.SEEDPROM
M0 5 221 9 5 N L=1.8e-07 W=1e-06 $X=156860 $Y=741655 $D=0
M1 5 515 471 5 N L=1.8e-07 W=4.2e-07 $X=325300 $Y=655750 $D=0
M2 678 82 5 5 N L=1.8e-07 W=4.2e-07 $X=326210 $Y=655750 $D=0
M3 515 516 678 5 N L=1.8e-07 W=4.2e-07 $X=326680 $Y=655750 $D=0
M4 221 221 4 4 P L=1.8e-07 W=1.37e-06 $X=156860 $Y=739425 $D=16
M5 4 515 471 4 P L=1.8e-07 W=1.13e-06 $X=325300 $Y=653370 $D=16
M6 515 82 4 4 P L=1.8e-07 W=7.55e-07 $X=325970 $Y=653745 $D=16
M7 4 516 515 4 P L=1.8e-07 W=7.1e-07 $X=326720 $Y=653790 $D=16
X19 3 4 5 5 2 9 384 6 9 677 9 5 PDDW0208CDG $T=0 690000 0 270 $X=0 $Y=609400
X180 4 5 DCAPBWP7T $T=156120 625400 0 0 $X=155830 $Y=625165
X181 4 5 DCAPBWP7T $T=156120 719480 1 0 $X=155830 $Y=715270
X182 4 5 DCAPBWP7T $T=156120 735160 1 0 $X=155830 $Y=730950
X183 4 5 DCAPBWP7T $T=160600 680280 0 0 $X=160310 $Y=680045
X184 4 5 DCAPBWP7T $T=162840 664600 1 0 $X=162550 $Y=660390
X185 4 5 DCAPBWP7T $T=165080 601880 0 0 $X=164790 $Y=601645
X186 4 5 DCAPBWP7T $T=167880 672440 0 0 $X=167590 $Y=672205
X187 4 5 DCAPBWP7T $T=174040 735160 0 0 $X=173750 $Y=734925
X188 4 5 DCAPBWP7T $T=178520 711640 1 0 $X=178230 $Y=707430
X189 4 5 DCAPBWP7T $T=178520 735160 1 0 $X=178230 $Y=730950
X190 4 5 DCAPBWP7T $T=195320 648920 0 0 $X=195030 $Y=648685
X191 4 5 DCAPBWP7T $T=195320 664600 1 0 $X=195030 $Y=660390
X192 4 5 DCAPBWP7T $T=237320 656760 1 0 $X=237030 $Y=652550
X193 4 5 DCAPBWP7T $T=240120 711640 1 0 $X=239830 $Y=707430
X194 4 5 DCAPBWP7T $T=249080 664600 0 0 $X=248790 $Y=664365
X195 4 5 DCAPBWP7T $T=291080 641080 1 0 $X=290790 $Y=636870
X196 4 5 DCAPBWP7T $T=321320 641080 0 0 $X=321030 $Y=640845
X197 4 5 DCAPBWP7T $T=321320 719480 1 0 $X=321030 $Y=715270
X198 4 5 DCAPBWP7T $T=333080 695960 1 0 $X=332790 $Y=691750
X199 4 5 DCAPBWP7T $T=335320 735160 0 0 $X=335030 $Y=734925
X200 4 5 DCAPBWP7T $T=343720 633240 0 0 $X=343430 $Y=633005
X201 4 5 DCAPBWP7T $T=363320 656760 1 0 $X=363030 $Y=652550
X202 4 5 DCAPBWP7T $T=363320 727320 0 0 $X=363030 $Y=727085
X203 4 5 DCAPBWP7T $T=375080 735160 1 0 $X=374790 $Y=730950
X204 4 5 DCAPBWP7T $T=379560 711640 0 0 $X=379270 $Y=711405
X205 4 5 DCAPBWP7T $T=382920 609720 1 0 $X=382630 $Y=605510
X206 4 5 DCAPBWP7T $T=405320 688120 1 0 $X=405030 $Y=683910
X207 4 5 DCAPBWP7T $T=408120 719480 0 0 $X=407830 $Y=719245
X208 4 5 DCAPBWP7T $T=417080 672440 1 0 $X=416790 $Y=668230
X209 4 5 DCAPBWP7T $T=421560 703800 1 0 $X=421270 $Y=699590
X210 4 5 DCAPBWP7T $T=425480 680280 0 0 $X=425190 $Y=680045
X211 4 5 DCAPBWP7T $T=435000 664600 0 0 $X=434710 $Y=664365
X212 4 5 DCAPBWP7T $T=447320 648920 1 0 $X=447030 $Y=644710
X213 4 5 DCAPBWP7T $T=447320 664600 0 0 $X=447030 $Y=664365
X214 4 5 DCAPBWP7T $T=447320 672440 0 0 $X=447030 $Y=672205
X215 5 4 DCAP8BWP7T $T=156120 680280 1 0 $X=155830 $Y=676070
X216 5 4 DCAP8BWP7T $T=156120 727320 0 0 $X=155830 $Y=727085
X217 5 4 DCAP8BWP7T $T=158360 617560 0 0 $X=158070 $Y=617325
X218 5 4 DCAP8BWP7T $T=174040 695960 0 0 $X=173750 $Y=695725
X219 5 4 DCAP8BWP7T $T=182440 735160 1 0 $X=182150 $Y=730950
X220 5 4 DCAP8BWP7T $T=191400 703800 1 0 $X=191110 $Y=699590
X221 5 4 DCAP8BWP7T $T=191960 633240 1 0 $X=191670 $Y=629030
X222 5 4 DCAP8BWP7T $T=191960 656760 0 0 $X=191670 $Y=656525
X223 5 4 DCAP8BWP7T $T=192520 648920 1 0 $X=192230 $Y=644710
X224 5 4 DCAP8BWP7T $T=192520 695960 0 0 $X=192230 $Y=695725
X225 5 4 DCAP8BWP7T $T=221640 680280 0 0 $X=221350 $Y=680045
X226 5 4 DCAP8BWP7T $T=233400 735160 1 0 $X=233110 $Y=730950
X227 5 4 DCAP8BWP7T $T=233960 633240 0 0 $X=233670 $Y=633005
X228 5 4 DCAP8BWP7T $T=233960 688120 0 0 $X=233670 $Y=687885
X229 5 4 DCAP8BWP7T $T=233960 727320 1 0 $X=233670 $Y=723110
X230 5 4 DCAP8BWP7T $T=234520 648920 0 0 $X=234230 $Y=648685
X231 5 4 DCAP8BWP7T $T=275960 625400 0 0 $X=275670 $Y=625165
X232 5 4 DCAP8BWP7T $T=275960 633240 1 0 $X=275670 $Y=629030
X233 5 4 DCAP8BWP7T $T=275960 695960 0 0 $X=275670 $Y=695725
X234 5 4 DCAP8BWP7T $T=275960 703800 0 0 $X=275670 $Y=703565
X235 5 4 DCAP8BWP7T $T=275960 727320 0 0 $X=275670 $Y=727085
X236 5 4 DCAP8BWP7T $T=275960 735160 0 0 $X=275670 $Y=734925
X237 5 4 DCAP8BWP7T $T=276520 609720 1 0 $X=276230 $Y=605510
X238 5 4 DCAP8BWP7T $T=276520 625400 1 0 $X=276230 $Y=621190
X239 5 4 DCAP8BWP7T $T=306760 735160 1 0 $X=306470 $Y=730950
X240 5 4 DCAP8BWP7T $T=317960 617560 0 0 $X=317670 $Y=617325
X241 5 4 DCAP8BWP7T $T=317960 664600 1 0 $X=317670 $Y=660390
X242 5 4 DCAP8BWP7T $T=318520 609720 1 0 $X=318230 $Y=605510
X243 5 4 DCAP8BWP7T $T=318520 625400 1 0 $X=318230 $Y=621190
X244 5 4 DCAP8BWP7T $T=318520 711640 1 0 $X=318230 $Y=707430
X245 5 4 DCAP8BWP7T $T=324120 727320 1 0 $X=323830 $Y=723110
X246 5 4 DCAP8BWP7T $T=359960 688120 1 0 $X=359670 $Y=683910
X247 5 4 DCAP8BWP7T $T=359960 727320 1 0 $X=359670 $Y=723110
X248 5 4 DCAP8BWP7T $T=360520 609720 1 0 $X=360230 $Y=605510
X249 5 4 DCAP8BWP7T $T=360520 641080 0 0 $X=360230 $Y=640845
X250 5 4 DCAP8BWP7T $T=360520 735160 0 0 $X=360230 $Y=734925
X251 5 4 DCAP8BWP7T $T=366120 609720 0 0 $X=365830 $Y=609485
X252 5 4 DCAP8BWP7T $T=366120 625400 0 0 $X=365830 $Y=625165
X253 5 4 DCAP8BWP7T $T=366120 633240 0 0 $X=365830 $Y=633005
X254 5 4 DCAP8BWP7T $T=401400 625400 0 0 $X=401110 $Y=625165
X255 5 4 DCAP8BWP7T $T=401400 656760 1 0 $X=401110 $Y=652550
X256 5 4 DCAP8BWP7T $T=401960 625400 1 0 $X=401670 $Y=621190
X257 5 4 DCAP8BWP7T $T=401960 672440 1 0 $X=401670 $Y=668230
X258 5 4 DCAP8BWP7T $T=401960 680280 1 0 $X=401670 $Y=676070
X259 5 4 DCAP8BWP7T $T=401960 680280 0 0 $X=401670 $Y=680045
X260 5 4 DCAP8BWP7T $T=401960 711640 1 0 $X=401670 $Y=707430
X261 5 4 DCAP8BWP7T $T=402520 601880 0 0 $X=402230 $Y=601645
X262 5 4 DCAP8BWP7T $T=402520 609720 1 0 $X=402230 $Y=605510
X263 5 4 DCAP8BWP7T $T=402520 617560 1 0 $X=402230 $Y=613350
X264 5 4 DCAP8BWP7T $T=402520 664600 0 0 $X=402230 $Y=664365
X265 5 4 DCAP8BWP7T $T=444520 601880 1 0 $X=444230 $Y=597670
X266 5 4 DCAP8BWP7T $T=444520 609720 1 0 $X=444230 $Y=605510
X267 5 4 DCAP8BWP7T $T=444520 641080 1 0 $X=444230 $Y=636870
X268 5 4 DCAP8BWP7T $T=444520 672440 1 0 $X=444230 $Y=668230
X269 5 4 DCAP8BWP7T $T=444520 680280 0 0 $X=444230 $Y=680045
X270 5 4 DCAP4BWP7T $T=156120 656760 1 0 $X=155830 $Y=652550
X271 5 4 DCAP4BWP7T $T=170680 727320 1 0 $X=170390 $Y=723110
X272 5 4 DCAP4BWP7T $T=181880 609720 1 0 $X=181590 $Y=605510
X273 5 4 DCAP4BWP7T $T=194200 664600 0 0 $X=193910 $Y=664365
X274 5 4 DCAP4BWP7T $T=198120 695960 1 0 $X=197830 $Y=691750
X275 5 4 DCAP4BWP7T $T=198120 703800 0 0 $X=197830 $Y=703565
X276 5 4 DCAP4BWP7T $T=213240 703800 0 0 $X=212950 $Y=703565
X277 5 4 DCAP4BWP7T $T=236760 625400 0 0 $X=236470 $Y=625165
X278 5 4 DCAP4BWP7T $T=278200 664600 1 0 $X=277910 $Y=660390
X279 5 4 DCAP4BWP7T $T=278200 672440 0 0 $X=277910 $Y=672205
X280 5 4 DCAP4BWP7T $T=282120 711640 1 0 $X=281830 $Y=707430
X281 5 4 DCAP4BWP7T $T=291080 609720 0 0 $X=290790 $Y=609485
X282 5 4 DCAP4BWP7T $T=303400 727320 1 0 $X=303110 $Y=723110
X283 5 4 DCAP4BWP7T $T=312360 695960 1 0 $X=312070 $Y=691750
X284 5 4 DCAP4BWP7T $T=320200 601880 0 0 $X=319910 $Y=601645
X285 5 4 DCAP4BWP7T $T=320200 617560 1 0 $X=319910 $Y=613350
X286 5 4 DCAP4BWP7T $T=320200 664600 0 0 $X=319910 $Y=664365
X287 5 4 DCAP4BWP7T $T=320760 656760 1 0 $X=320470 $Y=652550
X288 5 4 DCAP4BWP7T $T=324120 617560 1 0 $X=323830 $Y=613350
X289 5 4 DCAP4BWP7T $T=324120 648920 1 0 $X=323830 $Y=644710
X290 5 4 DCAP4BWP7T $T=366120 601880 1 0 $X=365830 $Y=597670
X291 5 4 DCAP4BWP7T $T=373400 672440 0 0 $X=373110 $Y=672205
X292 5 4 DCAP4BWP7T $T=377880 601880 1 0 $X=377590 $Y=597670
X293 5 4 DCAP4BWP7T $T=380120 648920 0 0 $X=379830 $Y=648685
X294 5 4 DCAP4BWP7T $T=404760 633240 0 0 $X=404470 $Y=633005
X295 5 4 DCAP4BWP7T $T=404760 711640 0 0 $X=404470 $Y=711405
X296 5 4 DCAP4BWP7T $T=408120 711640 0 0 $X=407830 $Y=711405
X297 5 4 DCAP4BWP7T $T=408120 727320 1 0 $X=407830 $Y=723110
X298 5 4 DCAP4BWP7T $T=408120 735160 0 0 $X=407830 $Y=734925
X299 5 4 DCAP4BWP7T $T=415400 680280 0 0 $X=415110 $Y=680045
X300 5 4 DCAP4BWP7T $T=417080 735160 1 0 $X=416790 $Y=730950
X301 5 4 DCAP4BWP7T $T=431640 641080 1 0 $X=431350 $Y=636870
X302 5 4 DCAP4BWP7T $T=435000 625400 0 0 $X=434710 $Y=625165
X303 5 4 DCAP4BWP7T $T=440040 672440 1 0 $X=439750 $Y=668230
X304 5 4 ICV_40 $T=156120 633240 0 0 $X=155830 $Y=633005
X305 5 4 ICV_40 $T=165080 688120 1 0 $X=164790 $Y=683910
X306 5 4 ICV_40 $T=173480 680280 0 0 $X=173190 $Y=680045
X307 5 4 ICV_40 $T=176280 719480 0 0 $X=175990 $Y=719245
X308 5 4 ICV_40 $T=179080 695960 1 0 $X=178790 $Y=691750
X309 5 4 ICV_40 $T=183000 688120 0 0 $X=182710 $Y=687885
X310 5 4 ICV_40 $T=189160 601880 1 0 $X=188870 $Y=597670
X311 5 4 ICV_40 $T=189160 641080 1 0 $X=188870 $Y=636870
X312 5 4 ICV_40 $T=189160 641080 0 0 $X=188870 $Y=640845
X313 5 4 ICV_40 $T=189160 672440 1 0 $X=188870 $Y=668230
X314 5 4 ICV_40 $T=189160 695960 1 0 $X=188870 $Y=691750
X315 5 4 ICV_40 $T=189160 735160 1 0 $X=188870 $Y=730950
X316 5 4 ICV_40 $T=189160 743000 1 0 $X=188870 $Y=738790
X317 5 4 ICV_40 $T=189720 609720 1 0 $X=189430 $Y=605510
X318 5 4 ICV_40 $T=189720 680280 1 0 $X=189430 $Y=676070
X319 5 4 ICV_40 $T=190280 617560 0 0 $X=189990 $Y=617325
X320 5 4 ICV_40 $T=190280 711640 0 0 $X=189990 $Y=711405
X321 5 4 ICV_40 $T=198120 672440 0 0 $X=197830 $Y=672205
X322 5 4 ICV_40 $T=207080 648920 0 0 $X=206790 $Y=648685
X323 5 4 ICV_40 $T=207080 656760 1 0 $X=206790 $Y=652550
X324 5 4 ICV_40 $T=207080 664600 0 0 $X=206790 $Y=664365
X325 5 4 ICV_40 $T=214920 680280 1 0 $X=214630 $Y=676070
X326 5 4 ICV_40 $T=220520 648920 1 0 $X=220230 $Y=644710
X327 5 4 ICV_40 $T=221640 743000 1 0 $X=221350 $Y=738790
X328 5 4 ICV_40 $T=225000 688120 1 0 $X=224710 $Y=683910
X329 5 4 ICV_40 $T=231160 664600 1 0 $X=230870 $Y=660390
X330 5 4 ICV_40 $T=231720 695960 1 0 $X=231430 $Y=691750
X331 5 4 ICV_40 $T=231720 743000 1 0 $X=231430 $Y=738790
X332 5 4 ICV_40 $T=232280 648920 1 0 $X=231990 $Y=644710
X333 5 4 ICV_40 $T=232280 680280 1 0 $X=231990 $Y=676070
X334 5 4 ICV_40 $T=249080 695960 0 0 $X=248790 $Y=695725
X335 5 4 ICV_40 $T=249640 633240 0 0 $X=249350 $Y=633005
X336 5 4 ICV_40 $T=273160 601880 1 0 $X=272870 $Y=597670
X337 5 4 ICV_40 $T=273160 735160 1 0 $X=272870 $Y=730950
X338 5 4 ICV_40 $T=273720 617560 1 0 $X=273430 $Y=613350
X339 5 4 ICV_40 $T=273720 680280 1 0 $X=273430 $Y=676070
X340 5 4 ICV_40 $T=273720 688120 1 0 $X=273430 $Y=683910
X341 5 4 ICV_40 $T=273720 727320 1 0 $X=273430 $Y=723110
X342 5 4 ICV_40 $T=274280 617560 0 0 $X=273990 $Y=617325
X343 5 4 ICV_40 $T=300040 617560 0 0 $X=299750 $Y=617325
X344 5 4 ICV_40 $T=302280 648920 0 0 $X=301990 $Y=648685
X345 5 4 ICV_40 $T=303960 625400 1 0 $X=303670 $Y=621190
X346 5 4 ICV_40 $T=307320 695960 0 0 $X=307030 $Y=695725
X347 5 4 ICV_40 $T=315160 633240 1 0 $X=314870 $Y=629030
X348 5 4 ICV_40 $T=316280 648920 1 0 $X=315990 $Y=644710
X349 5 4 ICV_40 $T=316280 735160 0 0 $X=315990 $Y=734925
X350 5 4 ICV_40 $T=324120 727320 0 0 $X=323830 $Y=727085
X351 5 4 ICV_40 $T=342040 609720 1 0 $X=341750 $Y=605510
X352 5 4 ICV_40 $T=358280 617560 1 0 $X=357990 $Y=613350
X353 5 4 ICV_40 $T=381800 625400 0 0 $X=381510 $Y=625165
X354 5 4 ICV_40 $T=385160 601880 1 0 $X=384870 $Y=597670
X355 5 4 ICV_40 $T=385160 641080 0 0 $X=384870 $Y=640845
X356 5 4 ICV_40 $T=400280 641080 1 0 $X=399990 $Y=636870
X357 5 4 ICV_40 $T=413160 711640 1 0 $X=412870 $Y=707430
X358 5 4 ICV_40 $T=420440 609720 0 0 $X=420150 $Y=609485
X359 5 4 ICV_40 $T=426040 625400 1 0 $X=425750 $Y=621190
X360 5 4 ICV_40 $T=426040 656760 1 0 $X=425750 $Y=652550
X361 5 4 ICV_40 $T=429400 641080 0 0 $X=429110 $Y=640845
X362 5 4 ICV_40 $T=429400 680280 0 0 $X=429110 $Y=680045
X363 5 4 ICV_40 $T=441160 735160 1 0 $X=440870 $Y=730950
X364 5 4 ICV_40 $T=441720 711640 0 0 $X=441430 $Y=711405
X365 5 4 ICV_40 $T=441720 727320 0 0 $X=441430 $Y=727085
X366 5 4 ICV_40 $T=442280 617560 1 0 $X=441990 $Y=613350
X367 5 4 ICV_40 $T=442280 633240 1 0 $X=441990 $Y=629030
X368 5 4 ICV_40 $T=442280 735160 0 0 $X=441990 $Y=734925
X369 10 4 222 12 5 NR2D1BWP7T $T=156120 617560 0 0 $X=155830 $Y=617325
X370 11 4 224 16 5 NR2D1BWP7T $T=157240 609720 1 0 $X=156950 $Y=605510
X371 12 4 229 16 5 NR2D1BWP7T $T=157800 625400 0 0 $X=157510 $Y=625165
X372 232 4 225 13 5 NR2D1BWP7T $T=160040 719480 0 180 $X=157510 $Y=715270
X373 17 4 233 15 5 NR2D1BWP7T $T=158360 656760 1 0 $X=158070 $Y=652550
X374 19 4 231 226 5 NR2D1BWP7T $T=161720 609720 0 180 $X=159190 $Y=605510
X375 10 4 241 226 5 NR2D1BWP7T $T=159480 648920 1 0 $X=159190 $Y=644710
X376 235 4 234 232 5 NR2D1BWP7T $T=161720 727320 0 180 $X=159190 $Y=723110
X377 20 4 227 18 5 NR2D1BWP7T $T=162280 601880 0 180 $X=159750 $Y=597670
X378 11 4 239 15 5 NR2D1BWP7T $T=160040 641080 1 0 $X=159750 $Y=636870
X379 235 4 242 246 5 NR2D1BWP7T $T=160600 727320 0 0 $X=160310 $Y=727085
X380 223 4 243 246 5 NR2D1BWP7T $T=160600 735160 1 0 $X=160310 $Y=730950
X381 11 4 245 10 5 NR2D1BWP7T $T=163960 609720 0 180 $X=161430 $Y=605510
X382 252 4 251 13 5 NR2D1BWP7T $T=165640 719480 0 180 $X=163110 $Y=715270
X383 246 4 250 13 5 NR2D1BWP7T $T=167880 719480 0 180 $X=165350 $Y=715270
X384 276 4 268 246 5 NR2D1BWP7T $T=175160 727320 0 180 $X=172630 $Y=723110
X385 258 4 272 13 5 NR2D1BWP7T $T=176280 719480 0 180 $X=173750 $Y=715270
X386 275 4 273 246 5 NR2D1BWP7T $T=176280 719480 1 180 $X=173750 $Y=719245
X387 30 4 279 13 5 NR2D1BWP7T $T=181320 719480 0 180 $X=178790 $Y=715270
X388 289 4 288 13 5 NR2D1BWP7T $T=182440 711640 0 180 $X=179910 $Y=707430
X389 289 4 291 285 5 NR2D1BWP7T $T=180200 735160 1 0 $X=179910 $Y=730950
X390 20 4 277 15 5 NR2D1BWP7T $T=185240 601880 1 180 $X=182710 $Y=601645
X391 17 4 32 16 5 NR2D1BWP7T $T=186360 609720 0 180 $X=183830 $Y=605510
X392 289 4 298 223 5 NR2D1BWP7T $T=186360 727320 0 180 $X=183830 $Y=723110
X393 275 4 299 252 5 NR2D1BWP7T $T=186920 719480 1 180 $X=184390 $Y=719245
X394 20 4 300 10 5 NR2D1BWP7T $T=187480 601880 1 180 $X=184950 $Y=601645
X395 18 4 301 17 5 NR2D1BWP7T $T=185240 633240 1 0 $X=184950 $Y=629030
X396 275 4 303 30 5 NR2D1BWP7T $T=185240 735160 0 0 $X=184950 $Y=734925
X397 276 4 308 252 5 NR2D1BWP7T $T=189160 735160 0 180 $X=186630 $Y=730950
X398 232 4 324 285 5 NR2D1BWP7T $T=200920 735160 1 180 $X=198390 $Y=734925
X399 232 4 332 223 5 NR2D1BWP7T $T=200920 735160 0 0 $X=200630 $Y=734925
X400 20 4 351 19 5 NR2D1BWP7T $T=213800 625400 0 180 $X=211270 $Y=621190
X401 276 4 352 232 5 NR2D1BWP7T $T=214360 735160 0 180 $X=211830 $Y=730950
X402 19 4 354 11 5 NR2D1BWP7T $T=215480 609720 1 180 $X=212950 $Y=609485
X403 30 4 358 276 5 NR2D1BWP7T $T=216600 735160 0 180 $X=214070 $Y=730950
X404 19 4 51 17 5 NR2D1BWP7T $T=215480 609720 0 0 $X=215190 $Y=609485
X405 17 4 350 21 5 NR2D1BWP7T $T=217720 609720 0 0 $X=217430 $Y=609485
X406 289 4 387 235 5 NR2D1BWP7T $T=229480 688120 0 0 $X=229190 $Y=687885
X407 276 4 390 258 5 NR2D1BWP7T $T=231720 688120 0 0 $X=231430 $Y=687885
X408 289 4 420 276 5 NR2D1BWP7T $T=259160 695960 1 180 $X=256630 $Y=695725
X409 275 4 441 289 5 NR2D1BWP7T $T=268680 695960 0 0 $X=268390 $Y=695725
X410 235 4 403 252 5 NR2D1BWP7T $T=283240 727320 1 0 $X=282950 $Y=723110
X411 463 4 455 13 5 NR2D1BWP7T $T=289400 664600 0 180 $X=286870 $Y=660390
X412 468 4 466 13 5 NR2D1BWP7T $T=295560 664600 1 180 $X=293030 $Y=664365
X413 477 4 469 13 5 NR2D1BWP7T $T=297800 664600 1 180 $X=295270 $Y=664365
X414 104 4 100 486 5 NR2D1BWP7T $T=306200 633240 0 180 $X=303670 $Y=629030
X415 498 4 487 468 5 NR2D1BWP7T $T=310680 656760 0 0 $X=310390 $Y=656525
X416 486 4 497 105 5 NR2D1BWP7T $T=314040 648920 1 0 $X=313750 $Y=644710
X417 486 4 508 468 5 NR2D1BWP7T $T=317960 664600 0 180 $X=315430 $Y=660390
X418 498 4 510 104 5 NR2D1BWP7T $T=318520 625400 0 180 $X=315990 $Y=621190
X419 486 4 513 106 5 NR2D1BWP7T $T=324680 672440 1 0 $X=324390 $Y=668230
X420 498 4 495 13 5 NR2D1BWP7T $T=326920 711640 0 180 $X=324390 $Y=707430
X421 498 4 519 463 5 NR2D1BWP7T $T=329160 664600 0 180 $X=326630 $Y=660390
X422 558 4 524 13 5 NR2D1BWP7T $T=330840 727320 0 180 $X=328310 $Y=723110
X423 528 4 527 105 5 NR2D1BWP7T $T=332520 711640 0 180 $X=329990 $Y=707430
X424 498 4 540 106 5 NR2D1BWP7T $T=336440 680280 0 0 $X=336150 $Y=680045
X425 543 4 545 106 5 NR2D1BWP7T $T=338120 703800 0 0 $X=337830 $Y=703565
X426 104 4 550 528 5 NR2D1BWP7T $T=340360 703800 0 0 $X=340070 $Y=703565
X427 543 4 559 463 5 NR2D1BWP7T $T=342600 703800 0 0 $X=342310 $Y=703565
X428 104 4 537 558 5 NR2D1BWP7T $T=344840 680280 1 0 $X=344550 $Y=676070
X429 558 4 562 463 5 NR2D1BWP7T $T=345400 680280 0 0 $X=345110 $Y=680045
X430 104 4 507 543 5 NR2D1BWP7T $T=349320 641080 0 0 $X=349030 $Y=640845
X431 543 4 544 468 5 NR2D1BWP7T $T=351000 680280 1 0 $X=350710 $Y=676070
X432 114 4 570 13 5 NR2D1BWP7T $T=354920 641080 1 180 $X=352390 $Y=640845
X433 543 4 582 105 5 NR2D1BWP7T $T=358280 641080 0 0 $X=357990 $Y=640845
X434 122 4 567 13 5 NR2D1BWP7T $T=368920 641080 1 180 $X=366390 $Y=640845
X435 477 4 588 486 5 NR2D1BWP7T $T=366680 656760 1 0 $X=366390 $Y=652550
X436 498 4 573 477 5 NR2D1BWP7T $T=366680 680280 1 0 $X=366390 $Y=676070
X437 104 4 533 592 5 NR2D1BWP7T $T=367240 703800 1 0 $X=366950 $Y=699590
X438 486 4 546 463 5 NR2D1BWP7T $T=371160 680280 0 180 $X=368630 $Y=676070
X439 124 4 125 126 5 NR2D1BWP7T $T=370040 601880 1 0 $X=369750 $Y=597670
X440 558 4 596 105 5 NR2D1BWP7T $T=372280 703800 1 180 $X=369750 $Y=703565
X441 127 4 131 611 5 NR2D1BWP7T $T=373960 641080 0 0 $X=373670 $Y=640845
X442 592 4 607 105 5 NR2D1BWP7T $T=375080 711640 0 0 $X=374790 $Y=711405
X443 127 4 129 124 5 NR2D1BWP7T $T=375640 601880 1 0 $X=375350 $Y=597670
X444 124 4 610 13 5 NR2D1BWP7T $T=378440 648920 1 0 $X=378150 $Y=644710
X445 130 4 132 133 5 NR2D1BWP7T $T=379560 625400 0 0 $X=379270 $Y=625165
X446 115 4 134 611 5 NR2D1BWP7T $T=380120 641080 1 0 $X=379830 $Y=636870
X447 468 4 566 592 5 NR2D1BWP7T $T=383480 711640 1 180 $X=380950 $Y=711405
X448 638 4 637 13 5 NR2D1BWP7T $T=392440 648920 0 0 $X=392150 $Y=648685
X449 611 4 639 139 5 NR2D1BWP7T $T=395240 601880 1 0 $X=394950 $Y=597670
X450 115 4 143 638 5 NR2D1BWP7T $T=400280 601880 0 0 $X=399990 $Y=601645
X451 638 4 656 139 5 NR2D1BWP7T $T=402520 609720 0 180 $X=399990 $Y=605510
X452 611 4 614 13 5 NR2D1BWP7T $T=410920 633240 0 180 $X=408390 $Y=629030
X453 486 4 506 13 5 NR2D1BWP7T $T=412600 727320 0 180 $X=410070 $Y=723110
X454 468 4 606 558 5 NR2D1BWP7T $T=410920 711640 1 0 $X=410630 $Y=707430
X455 543 4 505 13 5 NR2D1BWP7T $T=413720 719480 1 180 $X=411190 $Y=719245
X456 592 4 555 13 5 NR2D1BWP7T $T=414840 727320 1 180 $X=412310 $Y=727085
X457 149 4 648 13 5 NR2D1BWP7T $T=417640 735160 1 180 $X=415110 $Y=734925
X458 160 4 623 13 5 NR2D1BWP7T $T=421560 735160 0 180 $X=419030 $Y=730950
X459 153 4 574 13 5 NR2D1BWP7T $T=423240 727320 0 180 $X=420710 $Y=723110
X460 154 4 575 13 5 NR2D1BWP7T $T=423240 735160 1 180 $X=420710 $Y=734925
X461 528 4 490 13 5 NR2D1BWP7T $T=423800 711640 1 180 $X=421270 $Y=711405
X462 158 4 599 13 5 NR2D1BWP7T $T=425480 727320 0 180 $X=422950 $Y=723110
X463 159 4 625 13 5 NR2D1BWP7T $T=426040 735160 1 180 $X=423510 $Y=734925
X464 165 4 665 159 5 NR2D1BWP7T $T=425480 695960 0 0 $X=425190 $Y=695725
X465 154 4 166 164 5 NR2D1BWP7T $T=428280 688120 1 180 $X=425750 $Y=687885
X466 168 4 600 13 5 NR2D1BWP7T $T=428280 735160 1 180 $X=425750 $Y=734925
X467 164 4 171 168 5 NR2D1BWP7T $T=429400 680280 1 180 $X=426870 $Y=680045
X468 165 4 671 160 5 NR2D1BWP7T $T=429960 735160 1 0 $X=429670 $Y=730950
X469 154 4 180 181 5 NR2D1BWP7T $T=431640 735160 0 0 $X=431350 $Y=734925
X470 164 4 670 159 5 NR2D1BWP7T $T=434440 727320 0 180 $X=431910 $Y=723110
X471 159 4 185 181 5 NR2D1BWP7T $T=435000 735160 0 0 $X=434710 $Y=734925
X472 154 4 673 192 5 NR2D1BWP7T $T=436120 727320 1 0 $X=435830 $Y=723110
X473 198 4 676 189 5 NR2D1BWP7T $T=440600 664600 0 180 $X=438070 $Y=660390
X474 214 4 210 189 5 NR2D1BWP7T $T=444520 609720 0 180 $X=441990 $Y=605510
X475 215 4 209 207 5 NR2D1BWP7T $T=444520 672440 0 180 $X=441990 $Y=668230
X476 4 5 DCAP64BWP7T $T=157800 617560 1 0 $X=157510 $Y=613350
X477 4 5 DCAP64BWP7T $T=328040 719480 0 0 $X=327750 $Y=719245
X478 4 5 DCAP64BWP7T $T=329160 664600 1 0 $X=328870 $Y=660390
X479 4 5 DCAP64BWP7T $T=408120 633240 0 0 $X=407830 $Y=633005
X480 4 5 DCAP64BWP7T $T=408120 648920 0 0 $X=407830 $Y=648685
X481 4 5 DCAP64BWP7T $T=408120 695960 1 0 $X=407830 $Y=691750
X482 4 5 DCAP64BWP7T $T=408120 703800 0 0 $X=407830 $Y=703565
X483 4 5 DCAP64BWP7T $T=408120 719480 1 0 $X=407830 $Y=715270
X484 4 5 DCAP64BWP7T $T=408120 743000 1 0 $X=407830 $Y=738790
X485 5 4 ICV_46 $T=156120 609720 0 0 $X=155830 $Y=609485
X486 5 4 ICV_46 $T=198120 711640 1 0 $X=197830 $Y=707430
X487 5 4 ICV_46 $T=198120 711640 0 0 $X=197830 $Y=711405
X488 5 4 ICV_46 $T=240120 672440 1 0 $X=239830 $Y=668230
X489 5 4 ICV_46 $T=240120 703800 1 0 $X=239830 $Y=699590
X490 5 4 ICV_46 $T=282120 688120 0 0 $X=281830 $Y=687885
X491 5 4 ICV_46 $T=366120 727320 0 0 $X=365830 $Y=727085
X529 5 4 ICV_47 $T=156120 625400 1 0 $X=155830 $Y=621190
X530 5 4 ICV_47 $T=198120 641080 0 0 $X=197830 $Y=640845
X531 5 4 ICV_47 $T=198120 656760 0 0 $X=197830 $Y=656525
X532 5 4 ICV_47 $T=198120 672440 1 0 $X=197830 $Y=668230
X533 5 4 ICV_47 $T=240120 641080 0 0 $X=239830 $Y=640845
X534 5 4 ICV_47 $T=240120 711640 0 0 $X=239830 $Y=711405
X535 5 4 ICV_47 $T=240120 719480 1 0 $X=239830 $Y=715270
X536 5 4 ICV_47 $T=240120 743000 1 0 $X=239830 $Y=738790
X537 5 4 ICV_47 $T=282120 703800 1 0 $X=281830 $Y=699590
X538 5 4 ICV_47 $T=282120 711640 0 0 $X=281830 $Y=711405
X539 5 4 ICV_47 $T=282120 727320 0 0 $X=281830 $Y=727085
X540 5 4 ICV_47 $T=324120 601880 0 0 $X=323830 $Y=601645
X541 5 4 ICV_47 $T=324120 641080 1 0 $X=323830 $Y=636870
X542 5 4 ICV_47 $T=324120 656760 0 0 $X=323830 $Y=656525
X543 5 4 ICV_47 $T=324120 672440 0 0 $X=323830 $Y=672205
X544 5 4 ICV_47 $T=324120 688120 0 0 $X=323830 $Y=687885
X545 5 4 ICV_47 $T=324120 703800 1 0 $X=323830 $Y=699590
X546 5 4 ICV_47 $T=324120 735160 1 0 $X=323830 $Y=730950
X547 5 4 ICV_47 $T=324120 743000 1 0 $X=323830 $Y=738790
X548 5 4 ICV_47 $T=366120 633240 1 0 $X=365830 $Y=629030
X549 5 4 ICV_47 $T=366120 695960 1 0 $X=365830 $Y=691750
X550 5 4 ICV_47 $T=366120 743000 1 0 $X=365830 $Y=738790
X551 4 5 DCAP32BWP7T $T=166760 633240 1 0 $X=166470 $Y=629030
X552 4 5 DCAP32BWP7T $T=166760 703800 0 0 $X=166470 $Y=703565
X553 4 5 DCAP32BWP7T $T=177400 664600 1 0 $X=177110 $Y=660390
X554 4 5 DCAP32BWP7T $T=214920 617560 1 0 $X=214630 $Y=613350
X555 4 5 DCAP32BWP7T $T=221080 601880 1 0 $X=220790 $Y=597670
X556 4 5 DCAP32BWP7T $T=240120 656760 0 0 $X=239830 $Y=656525
X557 4 5 DCAP32BWP7T $T=240120 735160 1 0 $X=239830 $Y=730950
X558 4 5 DCAP32BWP7T $T=255800 617560 1 0 $X=255510 $Y=613350
X559 4 5 DCAP32BWP7T $T=258040 625400 0 0 $X=257750 $Y=625165
X560 4 5 DCAP32BWP7T $T=259160 680280 0 0 $X=258870 $Y=680045
X561 4 5 DCAP32BWP7T $T=262520 695960 1 0 $X=262230 $Y=691750
X562 4 5 DCAP32BWP7T $T=282120 648920 1 0 $X=281830 $Y=644710
X563 4 5 DCAP32BWP7T $T=282120 719480 1 0 $X=281830 $Y=715270
X564 4 5 DCAP32BWP7T $T=285480 727320 1 0 $X=285190 $Y=723110
X565 4 5 DCAP32BWP7T $T=300600 719480 0 0 $X=300310 $Y=719245
X566 4 5 DCAP32BWP7T $T=303960 609720 0 0 $X=303670 $Y=609485
X567 4 5 DCAP32BWP7T $T=304520 601880 1 0 $X=304230 $Y=597670
X568 4 5 DCAP32BWP7T $T=345400 656760 1 0 $X=345110 $Y=652550
X569 4 5 DCAP32BWP7T $T=345400 727320 0 0 $X=345110 $Y=727085
X570 4 5 DCAP32BWP7T $T=366120 656760 0 0 $X=365830 $Y=656525
X571 4 5 DCAP32BWP7T $T=371160 680280 1 0 $X=370870 $Y=676070
X572 4 5 DCAP32BWP7T $T=380680 648920 1 0 $X=380390 $Y=644710
X573 4 5 DCAP32BWP7T $T=382360 641080 1 0 $X=382070 $Y=636870
X574 4 5 DCAP32BWP7T $T=385160 719480 1 0 $X=384870 $Y=715270
X575 4 5 DCAP32BWP7T $T=386840 711640 0 0 $X=386550 $Y=711405
X576 4 5 DCAP32BWP7T $T=388520 672440 0 0 $X=388230 $Y=672205
X577 4 5 DCAP32BWP7T $T=388520 727320 1 0 $X=388230 $Y=723110
X578 4 5 DCAP32BWP7T $T=389080 703800 1 0 $X=388790 $Y=699590
X579 4 5 DCAP32BWP7T $T=408120 625400 1 0 $X=407830 $Y=621190
X580 4 5 DCAP32BWP7T $T=408120 656760 1 0 $X=407830 $Y=652550
X581 4 5 DCAP32BWP7T $T=408120 680280 1 0 $X=407830 $Y=676070
X582 4 5 DCAP32BWP7T $T=411480 641080 0 0 $X=411190 $Y=640845
X583 4 5 DCAP32BWP7T $T=424920 711640 1 0 $X=424630 $Y=707430
X584 4 5 DCAP32BWP7T $T=427720 703800 1 0 $X=427430 $Y=699590
X585 4 5 DCAP32BWP7T $T=430520 617560 0 0 $X=430230 $Y=617325
X586 229 241 239 269 4 5 274 FA1D0BWP7T $T=162840 617560 0 0 $X=162550 $Y=617325
X587 231 245 277 28 4 5 280 FA1D0BWP7T $T=166760 601880 0 0 $X=166470 $Y=601645
X588 278 233 227 259 4 5 255 FA1D0BWP7T $T=179640 648920 0 180 $X=166470 $Y=644710
X589 265 259 280 290 4 5 293 FA1D0BWP7T $T=170120 633240 0 0 $X=169830 $Y=633005
X590 247 224 222 313 4 5 316 FA1D0BWP7T $T=177400 617560 0 0 $X=177110 $Y=617325
X591 255 253 281 318 4 5 284 FA1D0BWP7T $T=179080 656760 0 0 $X=178790 $Y=656525
X592 290 313 38 39 4 5 41 FA1D0BWP7T $T=198680 601880 0 0 $X=198390 $Y=601645
X593 269 316 327 333 4 5 372 FA1D0BWP7T $T=198680 617560 0 0 $X=198390 $Y=617325
X594 318 333 293 40 4 5 346 FA1D0BWP7T $T=198680 633240 1 0 $X=198390 $Y=629030
X595 301 340 330 327 4 5 325 FA1D0BWP7T $T=211560 648920 0 180 $X=198390 $Y=644710
X596 291 234 299 328 4 5 326 FA1D0BWP7T $T=211560 719480 1 180 $X=198390 $Y=719245
X597 329 323 347 348 4 5 317 FA1D0BWP7T $T=200360 695960 1 0 $X=200070 $Y=691750
X598 328 336 345 347 4 5 304 FA1D0BWP7T $T=200360 703800 0 0 $X=200070 $Y=703565
X599 344 350 354 53 4 5 55 FA1D0BWP7T $T=208200 601880 1 0 $X=207910 $Y=597670
X600 309 257 268 345 4 5 349 FA1D0BWP7T $T=224440 719480 1 180 $X=211270 $Y=719245
X601 263 242 332 389 4 5 391 FA1D0BWP7T $T=220520 735160 1 0 $X=220230 $Y=730950
X602 352 298 273 376 4 5 336 FA1D0BWP7T $T=234520 719480 0 180 $X=221350 $Y=715270
X603 243 324 403 407 4 5 412 FA1D0BWP7T $T=240680 719480 0 0 $X=240390 $Y=719245
X604 343 400 326 408 4 5 413 FA1D0BWP7T $T=240680 735160 0 0 $X=240390 $Y=734925
X605 358 365 405 410 4 5 414 FA1D0BWP7T $T=241240 695960 1 0 $X=240950 $Y=691750
X606 408 389 349 315 4 5 395 FA1D0BWP7T $T=254680 711640 0 180 $X=241510 $Y=707430
X607 375 376 322 338 4 5 329 FA1D0BWP7T $T=263640 664600 1 180 $X=250470 $Y=664365
X608 409 334 426 431 4 5 433 FA1D0BWP7T $T=251880 727320 1 0 $X=251590 $Y=723110
X609 382 308 303 400 4 5 409 FA1D0BWP7T $T=266440 735160 1 180 $X=253270 $Y=734925
X610 407 391 410 437 4 5 439 FA1D0BWP7T $T=255800 711640 1 0 $X=255510 $Y=707430
X611 445 390 387 392 4 5 331 FA1D0BWP7T $T=273720 680280 0 180 $X=260550 $Y=676070
X612 425 424 394 434 4 5 406 FA1D0BWP7T $T=276520 664600 1 180 $X=263350 $Y=664365
X613 431 437 413 435 4 5 432 FA1D0BWP7T $T=276520 719480 1 180 $X=263350 $Y=719245
X614 363 435 395 501 4 5 503 FA1D0BWP7T $T=301720 672440 1 0 $X=301430 $Y=668230
X615 488 497 507 511 4 5 512 FA1D0BWP7T $T=305640 633240 0 0 $X=305350 $Y=633005
X616 494 107 518 534 4 5 538 FA1D0BWP7T $T=324680 601880 1 0 $X=324390 $Y=597670
X617 499 520 531 535 4 5 539 FA1D0BWP7T $T=324680 625400 0 0 $X=324390 $Y=625165
X618 525 532 546 549 4 5 552 FA1D0BWP7T $T=330280 664600 0 0 $X=329990 $Y=664365
X619 508 537 519 520 4 5 557 FA1D0BWP7T $T=332520 656760 1 0 $X=332230 $Y=652550
X620 533 544 540 554 4 5 563 FA1D0BWP7T $T=334760 695960 1 0 $X=334470 $Y=691750
X621 554 557 549 572 4 5 578 FA1D0BWP7T $T=343720 664600 0 0 $X=343430 $Y=664365
X622 539 565 572 576 4 5 579 FA1D0BWP7T $T=345960 648920 0 0 $X=345670 $Y=648685
X623 550 513 573 577 4 5 580 FA1D0BWP7T $T=345960 703800 0 0 $X=345670 $Y=703565
X624 562 566 545 581 4 5 584 FA1D0BWP7T $T=347640 695960 1 0 $X=347350 $Y=691750
X625 586 559 606 612 4 5 616 FA1D0BWP7T $T=366680 688120 0 0 $X=366390 $Y=687885
X626 588 603 618 620 4 5 622 FA1D0BWP7T $T=371160 664600 1 0 $X=370870 $Y=660390
X627 604 612 552 601 4 5 628 FA1D0BWP7T $T=375640 672440 0 0 $X=375350 $Y=672205
X628 605 577 563 604 4 5 631 FA1D0BWP7T $T=376200 703800 1 0 $X=375910 $Y=699590
X629 581 616 620 635 4 5 633 FA1D0BWP7T $T=379000 688120 1 0 $X=378710 $Y=683910
X630 608 640 628 627 4 5 624 FA1D0BWP7T $T=397480 609720 0 180 $X=384310 $Y=605510
X631 580 644 653 655 4 5 657 FA1D0BWP7T $T=389640 719480 0 0 $X=389350 $Y=719245
X632 655 635 631 640 4 5 652 FA1D0BWP7T $T=408680 695960 0 0 $X=408390 $Y=695725
X633 146 645 661 155 4 5 157 FA1D0BWP7T $T=412040 601880 1 0 $X=411750 $Y=597670
X634 670 673 671 674 4 5 204 FA1D0BWP7T $T=428840 711640 0 0 $X=428550 $Y=711405
X635 666 674 668 208 4 5 212 FA1D0BWP7T $T=431080 695960 0 0 $X=430790 $Y=695725
X636 7 5 4 12 INVD1BWP7T $T=156120 617560 1 0 $X=155830 $Y=613350
X637 14 5 4 11 INVD1BWP7T $T=158360 664600 1 180 $X=156390 $Y=664365
X638 220 5 4 15 INVD1BWP7T $T=156680 680280 0 0 $X=156390 $Y=680045
X639 228 5 4 223 INVD1BWP7T $T=159480 735160 0 180 $X=157510 $Y=730950
X640 218 5 4 16 INVD1BWP7T $T=159480 672440 1 0 $X=159190 $Y=668230
X641 249 5 4 10 INVD1BWP7T $T=173480 688120 0 180 $X=171510 $Y=683910
X642 27 5 4 246 INVD1BWP7T $T=177400 735160 1 180 $X=175430 $Y=734925
X643 295 5 4 276 INVD1BWP7T $T=183560 735160 1 180 $X=181590 $Y=734925
X644 314 5 4 19 INVD1BWP7T $T=191960 633240 0 180 $X=189990 $Y=629030
X645 362 5 4 355 INVD1BWP7T $T=223320 680280 0 180 $X=221350 $Y=676070
X646 442 5 4 232 INVD1BWP7T $T=270920 735160 1 180 $X=268950 $Y=734925
X647 369 5 4 289 INVD1BWP7T $T=272600 695960 1 180 $X=270630 $Y=695725
X648 448 5 4 252 INVD1BWP7T $T=273160 735160 0 180 $X=271190 $Y=730950
X649 450 5 4 460 INVD1BWP7T $T=287720 695960 0 0 $X=287430 $Y=695725
X650 514 5 4 468 INVD1BWP7T $T=348760 680280 0 180 $X=346790 $Y=676070
X651 595 5 4 558 INVD1BWP7T $T=385160 719480 0 180 $X=383190 $Y=715270
X652 140 5 4 611 INVD1BWP7T $T=398600 648920 1 180 $X=396630 $Y=648685
X653 142 5 4 141 INVD1BWP7T $T=401400 656760 0 180 $X=399430 $Y=652550
X654 594 5 4 592 INVD1BWP7T $T=411480 719480 1 180 $X=409510 $Y=719245
X655 663 5 4 463 INVD1BWP7T $T=419320 680280 1 180 $X=417350 $Y=680045
X656 646 5 4 477 INVD1BWP7T $T=426040 688120 1 180 $X=424070 $Y=687885
X657 598 5 4 106 INVD1BWP7T $T=427720 703800 0 180 $X=425750 $Y=699590
X658 379 5 4 667 INVD1BWP7T $T=426600 680280 1 0 $X=426310 $Y=676070
X659 197 5 4 175 INVD1BWP7T $T=440600 617560 1 0 $X=440310 $Y=613350
X795 7 5 237 240 4 ND2D1BWP7T $T=160040 641080 0 0 $X=159750 $Y=640845
X796 8 5 238 218 4 ND2D1BWP7T $T=160600 680280 1 0 $X=160310 $Y=676070
X797 7 5 244 220 4 ND2D1BWP7T $T=163400 672440 0 180 $X=160870 $Y=668230
X798 22 5 248 24 4 ND2D1BWP7T $T=162840 633240 0 0 $X=162550 $Y=633005
X799 228 5 260 261 4 ND2D1BWP7T $T=171240 743000 0 180 $X=168710 $Y=738790
X800 270 5 26 266 4 ND2D1BWP7T $T=174600 672440 1 180 $X=172070 $Y=672205
X801 8 5 264 240 4 ND2D1BWP7T $T=175720 688120 1 0 $X=175430 $Y=683910
X802 249 5 267 29 4 ND2D1BWP7T $T=177960 672440 1 0 $X=177670 $Y=668230
X803 294 5 31 286 4 ND2D1BWP7T $T=183000 672440 1 180 $X=180470 $Y=672205
X804 310 5 305 240 4 ND2D1BWP7T $T=188600 672440 1 180 $X=186070 $Y=672205
X805 312 5 306 261 4 ND2D1BWP7T $T=188600 727320 0 180 $X=186070 $Y=723110
X806 14 5 44 240 4 ND2D1BWP7T $T=212680 617560 1 0 $X=212390 $Y=613350
X807 14 5 357 48 4 ND2D1BWP7T $T=217720 625400 0 180 $X=215190 $Y=621190
X808 364 5 361 42 4 ND2D1BWP7T $T=218840 648920 1 180 $X=216310 $Y=648685
X809 292 5 337 261 4 ND2D1BWP7T $T=221640 743000 0 180 $X=219110 $Y=738790
X810 42 5 359 240 4 ND2D1BWP7T $T=228360 633240 1 180 $X=225830 $Y=633005
X811 385 5 65 360 4 ND2D1BWP7T $T=230600 633240 1 180 $X=228070 $Y=633005
X812 380 5 67 319 4 ND2D1BWP7T $T=228360 664600 0 0 $X=228070 $Y=664365
X813 386 5 384 368 4 ND2D1BWP7T $T=231160 664600 0 180 $X=228630 $Y=660390
X814 402 5 383 314 4 ND2D1BWP7T $T=249640 625400 0 180 $X=247110 $Y=621190
X815 415 5 85 399 4 ND2D1BWP7T $T=255800 617560 0 180 $X=253270 $Y=613350
X816 442 5 449 388 4 ND2D1BWP7T $T=275960 735160 1 180 $X=273430 $Y=734925
X817 295 5 458 456 4 ND2D1BWP7T $T=290520 735160 1 180 $X=287990 $Y=734925
X818 228 5 483 448 4 ND2D1BWP7T $T=305640 719480 0 180 $X=303110 $Y=715270
X819 292 5 491 27 4 ND2D1BWP7T $T=307880 719480 0 180 $X=305350 $Y=715270
X820 479 5 447 261 4 ND2D1BWP7T $T=316840 695960 0 180 $X=314310 $Y=691750
X821 480 5 521 522 4 ND2D1BWP7T $T=327480 656760 1 0 $X=327190 $Y=652550
X822 473 5 526 479 4 ND2D1BWP7T $T=329720 680280 0 0 $X=329430 $Y=680045
X823 583 5 587 121 4 ND2D1BWP7T $T=366680 617560 0 0 $X=366390 $Y=617325
X824 560 5 589 646 4 ND2D1BWP7T $T=366680 664600 0 0 $X=366390 $Y=664365
X825 481 5 530 369 4 ND2D1BWP7T $T=366680 703800 0 0 $X=366390 $Y=703565
X826 514 5 590 591 4 ND2D1BWP7T $T=371160 672440 1 180 $X=368630 $Y=672205
X827 595 5 597 598 4 ND2D1BWP7T $T=371160 672440 0 0 $X=370870 $Y=672205
X828 135 5 621 480 4 ND2D1BWP7T $T=385160 601880 0 180 $X=382630 $Y=597670
X829 568 5 649 482 4 ND2D1BWP7T $T=402520 656760 1 180 $X=399990 $Y=656525
X830 516 5 643 522 4 ND2D1BWP7T $T=410920 711640 0 180 $X=408390 $Y=707430
X831 57 5 462 261 4 ND2D1BWP7T $T=410360 735160 0 0 $X=410070 $Y=734925
X832 312 5 551 564 4 ND2D1BWP7T $T=418200 727320 1 0 $X=417910 $Y=723110
X833 594 5 647 663 4 ND2D1BWP7T $T=419320 711640 0 0 $X=419030 $Y=711405
X834 161 5 672 178 4 ND2D1BWP7T $T=433880 672440 1 180 $X=431350 $Y=672205
X835 203 5 669 178 4 ND2D1BWP7T $T=440600 727320 0 180 $X=438070 $Y=723110
X855 8 5 4 226 INVD0BWP7T $T=156680 664600 1 0 $X=156390 $Y=660390
X856 256 5 4 254 INVD0BWP7T $T=166200 711640 0 0 $X=165910 $Y=711405
X857 283 5 4 236 INVD0BWP7T $T=179640 672440 1 180 $X=177670 $Y=672205
X858 292 5 4 285 INVD0BWP7T $T=181880 735160 1 180 $X=179910 $Y=734925
X859 302 5 4 307 INVD0BWP7T $T=186360 719480 1 0 $X=186070 $Y=715270
X860 321 5 4 323 INVD0BWP7T $T=190840 688120 0 0 $X=190550 $Y=687885
X861 46 5 4 230 INVD0BWP7T $T=215480 625400 0 180 $X=213510 $Y=621190
X862 353 5 4 342 INVD0BWP7T $T=213800 735160 0 0 $X=213510 $Y=734925
X863 429 5 4 375 INVD0BWP7T $T=223320 703800 1 180 $X=221350 $Y=703565
X864 392 5 4 394 INVD0BWP7T $T=232840 688120 1 0 $X=232550 $Y=683910
X865 73 5 4 72 INVD0BWP7T $T=242360 601880 1 180 $X=240390 $Y=601645
X866 406 5 4 335 INVD0BWP7T $T=245720 641080 0 180 $X=243750 $Y=636870
X867 418 5 4 436 INVD0BWP7T $T=256920 641080 0 180 $X=254950 $Y=636870
X868 478 5 4 99 INVD0BWP7T $T=301160 633240 0 180 $X=299190 $Y=629030
X869 489 5 4 499 INVD0BWP7T $T=310120 656760 1 0 $X=309830 $Y=652550
X870 511 5 4 518 INVD0BWP7T $T=326360 617560 1 0 $X=326070 $Y=613350
X871 538 5 4 548 INVD0BWP7T $T=342040 617560 0 180 $X=340070 $Y=613350
X872 556 5 4 565 INVD0BWP7T $T=366680 648920 0 0 $X=366390 $Y=648685
X873 123 5 4 120 INVD0BWP7T $T=370040 601880 0 180 $X=368070 $Y=597670
X874 152 5 4 638 INVD0BWP7T $T=422680 641080 0 180 $X=420710 $Y=636870
X875 664 5 4 666 INVD0BWP7T $T=425480 719480 1 180 $X=423510 $Y=719245
X876 83 5 4 173 INVD0BWP7T $T=434440 727320 1 0 $X=434150 $Y=723110
X877 186 5 4 190 INVD0BWP7T $T=436680 664600 0 0 $X=436390 $Y=664365
X878 194 5 4 193 INVD0BWP7T $T=438920 625400 1 180 $X=436950 $Y=625165
X879 211 5 4 213 INVD0BWP7T $T=442840 601880 1 0 $X=442550 $Y=597670
X880 304 311 315 317 5 4 OAI21D0BWP7T $T=187480 711640 0 0 $X=187190 $Y=711405
X881 428 423 366 429 5 4 OAI21D0BWP7T $T=261400 695960 0 0 $X=261110 $Y=695725
X882 374 452 441 418 5 4 OAI21D0BWP7T $T=285480 680280 1 180 $X=282390 $Y=680045
X883 578 602 601 579 5 4 OAI21D0BWP7T $T=376200 648920 1 180 $X=373110 $Y=648685
X920 296 5 29 240 4 282 ND3D0BWP7T $T=184680 695960 1 180 $X=181590 $Y=695725
X921 36 5 42 249 4 33 ND3D0BWP7T $T=213240 609720 1 180 $X=210150 $Y=609485
X922 320 5 388 261 4 454 ND3D0BWP7T $T=285480 735160 0 0 $X=285190 $Y=734925
X923 467 5 480 482 4 478 ND3D0BWP7T $T=301160 633240 1 0 $X=300870 $Y=629030
X924 366 5 479 442 4 429 ND3D0BWP7T $T=306200 680280 1 0 $X=305910 $Y=676070
X925 485 5 480 514 4 489 ND3D0BWP7T $T=324680 664600 0 0 $X=324390 $Y=664365
X926 658 5 152 138 4 147 ND3D0BWP7T $T=420440 609720 1 180 $X=417350 $Y=609485
X927 541 5 591 522 4 636 ND3D0BWP7T $T=426040 703800 0 180 $X=422950 $Y=699590
X928 70 5 161 163 4 664 ND3D0BWP7T $T=424360 688120 1 0 $X=424070 $Y=683910
X929 5 4 DCAP16BWP7T $T=157800 743000 1 0 $X=157510 $Y=738790
X930 5 4 DCAP16BWP7T $T=161720 727320 1 0 $X=161430 $Y=723110
X931 5 4 DCAP16BWP7T $T=162840 727320 0 0 $X=162550 $Y=727085
X932 5 4 DCAP16BWP7T $T=169560 735160 1 0 $X=169270 $Y=730950
X933 5 4 DCAP16BWP7T $T=174040 688120 0 0 $X=173750 $Y=687885
X934 5 4 DCAP16BWP7T $T=175160 727320 1 0 $X=174870 $Y=723110
X935 5 4 DCAP16BWP7T $T=180200 641080 1 0 $X=179910 $Y=636870
X936 5 4 DCAP16BWP7T $T=186920 719480 0 0 $X=186630 $Y=719245
X937 5 4 DCAP16BWP7T $T=187480 601880 0 0 $X=187190 $Y=601645
X938 5 4 DCAP16BWP7T $T=198120 609720 0 0 $X=197830 $Y=609485
X939 5 4 DCAP16BWP7T $T=198120 625400 1 0 $X=197830 $Y=621190
X940 5 4 DCAP16BWP7T $T=198120 656760 1 0 $X=197830 $Y=652550
X941 5 4 DCAP16BWP7T $T=198120 664600 0 0 $X=197830 $Y=664365
X942 5 4 DCAP16BWP7T $T=211560 648920 1 0 $X=211270 $Y=644710
X943 5 4 DCAP16BWP7T $T=222760 695960 1 0 $X=222470 $Y=691750
X944 5 4 DCAP16BWP7T $T=223320 680280 1 0 $X=223030 $Y=676070
X945 5 4 DCAP16BWP7T $T=228920 601880 0 0 $X=228630 $Y=601645
X946 5 4 DCAP16BWP7T $T=229480 609720 1 0 $X=229190 $Y=605510
X947 5 4 DCAP16BWP7T $T=229480 609720 0 0 $X=229190 $Y=609485
X948 5 4 DCAP16BWP7T $T=229480 617560 0 0 $X=229190 $Y=617325
X949 5 4 DCAP16BWP7T $T=240120 727320 1 0 $X=239830 $Y=723110
X950 5 4 DCAP16BWP7T $T=244040 625400 0 0 $X=243750 $Y=625165
X951 5 4 DCAP16BWP7T $T=253560 625400 1 0 $X=253270 $Y=621190
X952 5 4 DCAP16BWP7T $T=253560 719480 0 0 $X=253270 $Y=719245
X953 5 4 DCAP16BWP7T $T=263640 609720 0 0 $X=263350 $Y=609485
X954 5 4 DCAP16BWP7T $T=264760 727320 1 0 $X=264470 $Y=723110
X955 5 4 DCAP16BWP7T $T=265320 617560 0 0 $X=265030 $Y=617325
X956 5 4 DCAP16BWP7T $T=269240 664600 1 0 $X=268950 $Y=660390
X957 5 4 DCAP16BWP7T $T=269240 672440 0 0 $X=268950 $Y=672205
X958 5 4 DCAP16BWP7T $T=270920 648920 1 0 $X=270630 $Y=644710
X959 5 4 DCAP16BWP7T $T=271480 656760 1 0 $X=271190 $Y=652550
X960 5 4 DCAP16BWP7T $T=272040 656760 0 0 $X=271750 $Y=656525
X961 5 4 DCAP16BWP7T $T=293320 648920 0 0 $X=293030 $Y=648685
X962 5 4 DCAP16BWP7T $T=296120 656760 1 0 $X=295830 $Y=652550
X963 5 4 DCAP16BWP7T $T=297240 711640 1 0 $X=296950 $Y=707430
X964 5 4 DCAP16BWP7T $T=307320 735160 0 0 $X=307030 $Y=734925
X965 5 4 DCAP16BWP7T $T=312920 656760 0 0 $X=312630 $Y=656525
X966 5 4 DCAP16BWP7T $T=312920 680280 0 0 $X=312630 $Y=680045
X967 5 4 DCAP16BWP7T $T=313480 641080 1 0 $X=313190 $Y=636870
X968 5 4 DCAP16BWP7T $T=313480 735160 1 0 $X=313190 $Y=730950
X969 5 4 DCAP16BWP7T $T=334200 727320 0 0 $X=333910 $Y=727085
X970 5 4 DCAP16BWP7T $T=342040 617560 1 0 $X=341750 $Y=613350
X971 5 4 DCAP16BWP7T $T=352120 609720 0 0 $X=351830 $Y=609485
X972 5 4 DCAP16BWP7T $T=354920 719480 1 0 $X=354630 $Y=715270
X973 5 4 DCAP16BWP7T $T=356040 633240 0 0 $X=355750 $Y=633005
X974 5 4 DCAP16BWP7T $T=366120 601880 0 0 $X=365830 $Y=601645
X975 5 4 DCAP16BWP7T $T=366120 641080 1 0 $X=365830 $Y=636870
X976 5 4 DCAP16BWP7T $T=366120 688120 1 0 $X=365830 $Y=683910
X977 5 4 DCAP16BWP7T $T=366120 727320 1 0 $X=365830 $Y=723110
X978 5 4 DCAP16BWP7T $T=366120 735160 1 0 $X=365830 $Y=730950
X979 5 4 DCAP16BWP7T $T=372280 703800 0 0 $X=371990 $Y=703565
X980 5 4 DCAP16BWP7T $T=377320 719480 0 0 $X=377030 $Y=719245
X981 5 4 DCAP16BWP7T $T=384040 617560 1 0 $X=383750 $Y=613350
X982 5 4 DCAP16BWP7T $T=394680 617560 0 0 $X=394390 $Y=617325
X983 5 4 DCAP16BWP7T $T=395800 633240 0 0 $X=395510 $Y=633005
X984 5 4 DCAP16BWP7T $T=397480 601880 1 0 $X=397190 $Y=597670
X985 5 4 DCAP16BWP7T $T=398040 664600 1 0 $X=397750 $Y=660390
X986 5 4 DCAP16BWP7T $T=408120 672440 1 0 $X=407830 $Y=668230
X987 5 4 DCAP16BWP7T $T=408120 735160 1 0 $X=407830 $Y=730950
X988 5 4 DCAP16BWP7T $T=413720 719480 0 0 $X=413430 $Y=719245
X989 5 4 DCAP16BWP7T $T=419320 672440 0 0 $X=419030 $Y=672205
X990 5 4 DCAP16BWP7T $T=422680 641080 1 0 $X=422390 $Y=636870
X991 5 4 DCAP16BWP7T $T=426040 664600 1 0 $X=425750 $Y=660390
X992 5 4 DCAP16BWP7T $T=426040 664600 0 0 $X=425750 $Y=664365
X993 5 4 DCAP16BWP7T $T=429960 609720 1 0 $X=429670 $Y=605510
X994 5 4 DCAP16BWP7T $T=431640 656760 0 0 $X=431350 $Y=656525
X995 5 4 DCAP16BWP7T $T=432200 735160 1 0 $X=431910 $Y=730950
X996 5 4 DCAP16BWP7T $T=433320 633240 1 0 $X=433030 $Y=629030
X997 5 4 DCAP16BWP7T $T=438360 664600 0 0 $X=438070 $Y=664365
X998 5 4 DCAP16BWP7T $T=438920 625400 0 0 $X=438630 $Y=625165
X1047 21 5 226 236 253 4 NR3D1BWP7T $T=159480 648920 0 0 $X=159190 $Y=648685
X1048 258 5 223 254 263 4 NR3D1BWP7T $T=172360 727320 0 0 $X=172070 $Y=727085
X1049 258 5 235 307 309 4 NR3D1BWP7T $T=192520 703800 1 180 $X=187750 $Y=703565
X1050 258 5 285 342 334 4 NR3D1BWP7T $T=213800 735160 1 180 $X=209030 $Y=734925
X1051 21 5 20 355 344 4 NR3D1BWP7T $T=245160 625400 0 180 $X=240390 $Y=621190
X1052 258 5 275 416 445 4 NR3D1BWP7T $T=274280 711640 0 180 $X=269510 $Y=707430
X1053 105 5 498 460 488 4 NR3D1BWP7T $T=338680 641080 0 0 $X=338390 $Y=640845
X1054 168 5 165 667 182 4 NR3D1BWP7T $T=432760 688120 1 0 $X=432470 $Y=683910
X1055 168 5 181 196 206 4 NR3D1BWP7T $T=437800 735160 0 0 $X=437510 $Y=734925
X1056 331 335 5 4 338 321 MAOI222D1BWP7T $T=201480 680280 1 0 $X=201190 $Y=676070
X1057 436 420 5 4 430 424 MAOI222D1BWP7T $T=265320 648920 1 180 $X=260550 $Y=648685
X1058 548 535 5 4 512 556 MAOI222D1BWP7T $T=345960 625400 0 180 $X=341190 $Y=621190
X1059 230 237 5 247 23 4 AOI21D1BWP7T $T=160600 633240 1 0 $X=160310 $Y=629030
X1060 254 260 5 263 257 4 AOI21D1BWP7T $T=166200 735160 1 0 $X=165910 $Y=730950
X1061 307 306 5 309 322 4 AOI21D1BWP7T $T=189160 695960 0 0 $X=188870 $Y=695725
X1062 342 337 5 334 343 4 AOI21D1BWP7T $T=206520 735160 1 180 $X=202870 $Y=734925
X1063 447 416 5 445 443 4 AOI21D1BWP7T $T=272600 695960 0 0 $X=272310 $Y=695725
X1064 447 416 5 445 430 4 AOI21D1BWP7T $T=286040 695960 1 180 $X=282390 $Y=695725
X1065 460 521 5 488 110 4 AOI21D1BWP7T $T=329160 641080 0 0 $X=328870 $Y=640845
X1066 175 170 5 659 172 4 AOI21D1BWP7T $T=429960 609720 0 180 $X=426310 $Y=605510
X1067 175 170 5 659 184 4 AOI21D1BWP7T $T=435560 601880 1 180 $X=431910 $Y=601645
X1068 240 21 4 5 INVD2BWP7T $T=165640 672440 0 0 $X=165350 $Y=672205
X1069 261 258 4 5 INVD2BWP7T $T=169000 743000 0 180 $X=166470 $Y=738790
X1070 370 416 4 5 INVD2BWP7T $T=253000 641080 1 0 $X=252710 $Y=636870
X1071 482 104 4 5 INVD2BWP7T $T=312920 625400 0 180 $X=310390 $Y=621190
X1072 479 275 4 5 INVD2BWP7T $T=315160 695960 0 0 $X=314870 $Y=695725
X1073 480 498 4 5 INVD2BWP7T $T=329160 641080 1 180 $X=326630 $Y=640845
X1074 312 235 4 5 INVD2BWP7T $T=345400 727320 1 180 $X=342870 $Y=727085
X1075 116 115 4 5 INVD2BWP7T $T=358280 617560 0 180 $X=355750 $Y=613350
X1076 522 105 4 5 INVD2BWP7T $T=357160 680280 1 0 $X=356870 $Y=676070
X1077 583 486 4 5 INVD2BWP7T $T=370600 648920 1 180 $X=368070 $Y=648685
X1078 199 205 4 5 INVD2BWP7T $T=440600 601880 1 0 $X=440310 $Y=597670
X1129 25 225 5 4 219 DFQD0BWP7T $T=166760 703800 1 180 $X=155830 $Y=703565
X1130 25 250 5 4 218 DFQD0BWP7T $T=167320 695960 0 180 $X=156390 $Y=691750
X1131 25 251 5 4 220 DFQD0BWP7T $T=168440 695960 1 0 $X=168150 $Y=691750
X1132 25 279 5 4 48 DFQD0BWP7T $T=204840 672440 0 0 $X=204550 $Y=672205
X1133 25 69 5 4 283 DFQD0BWP7T $T=234520 648920 1 180 $X=223590 $Y=648685
X1134 25 397 5 4 366 DFQD0BWP7T $T=240680 664600 1 0 $X=240390 $Y=660390
X1135 25 396 5 4 302 DFQD0BWP7T $T=240680 672440 0 0 $X=240390 $Y=672205
X1136 25 79 5 4 296 DFQD0BWP7T $T=254680 648920 0 180 $X=243750 $Y=644710
X1137 25 417 5 4 401 DFQD0BWP7T $T=259160 680280 1 180 $X=248230 $Y=680045
X1138 25 89 5 4 362 DFQD0BWP7T $T=265320 617560 1 180 $X=254390 $Y=617325
X1139 25 90 5 4 341 DFQD0BWP7T $T=267000 633240 1 180 $X=256070 $Y=633005
X1140 25 438 5 4 370 DFQD0BWP7T $T=270920 648920 0 180 $X=259990 $Y=644710
X1141 25 440 5 4 422 DFQD0BWP7T $T=272040 656760 1 180 $X=261110 $Y=656525
X1142 25 421 5 4 353 DFQD0BWP7T $T=273720 688120 0 180 $X=262790 $Y=683910
X1143 25 92 5 4 310 DFQD0BWP7T $T=276520 625400 0 180 $X=265590 $Y=621190
X1144 25 95 5 4 402 DFQD0BWP7T $T=293320 601880 1 180 $X=282390 $Y=601645
X1145 25 94 5 4 93 DFQD0BWP7T $T=293320 617560 0 180 $X=282390 $Y=613350
X1146 25 459 5 4 364 DFQD0BWP7T $T=293320 633240 0 180 $X=282390 $Y=629030
X1147 25 464 5 4 450 DFQD0BWP7T $T=295560 641080 1 180 $X=284630 $Y=640845
X1148 25 465 5 4 451 DFQD0BWP7T $T=295560 672440 0 180 $X=284630 $Y=668230
X1149 25 461 5 4 419 DFQD0BWP7T $T=296120 656760 0 180 $X=285190 $Y=652550
X1150 25 470 5 4 373 DFQD0BWP7T $T=298920 680280 1 180 $X=287990 $Y=680045
X1151 25 471 5 4 453 DFQD0BWP7T $T=298920 695960 0 180 $X=287990 $Y=691750
X1152 25 466 5 4 97 DFQD0BWP7T $T=303960 609720 1 180 $X=293030 $Y=609485
X1153 25 455 5 4 96 DFQD0BWP7T $T=303960 625400 0 180 $X=293030 $Y=621190
X1154 25 469 5 4 98 DFQD0BWP7T $T=304520 601880 0 180 $X=293590 $Y=597670
X1155 25 490 5 4 475 DFQD0BWP7T $T=309560 703800 1 180 $X=298630 $Y=703565
X1156 25 496 5 4 481 DFQD0BWP7T $T=312920 680280 1 180 $X=301990 $Y=680045
X1157 25 504 5 4 485 DFQD0BWP7T $T=317960 617560 1 180 $X=307030 $Y=617325
X1158 25 505 5 4 493 DFQD0BWP7T $T=318520 711640 0 180 $X=307590 $Y=707430
X1159 25 506 5 4 492 DFQD0BWP7T $T=318520 727320 0 180 $X=307590 $Y=723110
X1160 25 524 5 4 500 DFQD0BWP7T $T=335320 735160 1 180 $X=324390 $Y=734925
X1161 25 111 5 4 467 DFQD0BWP7T $T=340360 609720 1 180 $X=329430 $Y=609485
X1162 25 569 5 4 536 DFQD0BWP7T $T=356040 633240 1 180 $X=345110 $Y=633005
X1163 25 570 5 4 560 DFQD0BWP7T $T=356600 625400 0 180 $X=345670 $Y=621190
X1164 25 574 5 4 564 DFQD0BWP7T $T=359960 727320 0 180 $X=349030 $Y=723110
X1165 25 567 5 4 583 DFQD0BWP7T $T=349880 609720 1 0 $X=349590 $Y=605510
X1166 25 575 5 4 517 DFQD0BWP7T $T=360520 735160 1 180 $X=349590 $Y=734925
X1167 25 599 5 4 585 DFQD0BWP7T $T=377320 719480 1 180 $X=366390 $Y=719245
X1168 25 610 5 4 595 DFQD0BWP7T $T=381240 633240 1 180 $X=370310 $Y=633005
X1169 25 614 5 4 593 DFQD0BWP7T $T=381800 617560 1 180 $X=370870 $Y=617325
X1170 25 623 5 4 609 DFQD0BWP7T $T=387960 735160 1 180 $X=377030 $Y=734925
X1171 25 625 5 4 529 DFQD0BWP7T $T=388520 727320 0 180 $X=377590 $Y=723110
X1172 25 637 5 4 619 DFQD0BWP7T $T=394680 617560 1 180 $X=383750 $Y=617325
X1173 25 615 5 4 626 DFQD0BWP7T $T=395800 633240 1 180 $X=384870 $Y=633005
X1174 25 648 5 4 632 DFQD0BWP7T $T=400840 735160 1 180 $X=389910 $Y=734925
X1175 25 654 5 4 571 DFQD0BWP7T $T=419880 656760 1 180 $X=408950 $Y=656525
X1176 150 662 5 4 660 DFQD0BWP7T $T=421560 633240 0 180 $X=410630 $Y=629030
X1177 25 174 5 4 663 DFQD0BWP7T $T=431640 656760 1 180 $X=420710 $Y=656525
X1178 150 177 5 4 598 DFQD0BWP7T $T=433880 648920 0 180 $X=422950 $Y=644710
X1179 150 183 5 4 136 DFQD0BWP7T $T=438360 609720 1 180 $X=427430 $Y=609485
X1180 150 676 5 4 646 DFQD0BWP7T $T=444520 641080 0 180 $X=433590 $Y=636870
X1181 230 5 4 12 21 247 NR3D0BWP7T $T=163960 633240 1 0 $X=163670 $Y=629030
X1182 344 4 47 359 355 5 AOI21D2BWP7T $T=218840 625400 1 180 $X=213510 $Y=625165
X1183 182 4 187 672 667 5 AOI21D2BWP7T $T=440040 672440 0 180 $X=434710 $Y=668230
X1184 264 265 236 253 5 4 AOI21D0BWP7T $T=169560 672440 0 0 $X=169270 $Y=672205
X1185 521 484 460 488 5 4 AOI21D0BWP7T $T=329160 648920 0 180 $X=326070 $Y=644710
X1186 669 668 173 169 5 4 AOI21D0BWP7T $T=429960 727320 0 180 $X=426870 $Y=723110
X1187 356 5 4 360 BUFFD0BWP7T $T=213800 656760 1 0 $X=213510 $Y=652550
X1188 423 5 4 425 BUFFD0BWP7T $T=259160 695960 0 0 $X=258870 $Y=695725
X1189 29 240 5 4 287 AN2D1BWP7T $T=189160 695960 0 180 $X=186070 $Y=691750
X1190 29 314 5 4 278 AN2D1BWP7T $T=190280 633240 0 180 $X=187190 $Y=629030
X1191 24 42 5 4 330 AN2D1BWP7T $T=216600 648920 1 180 $X=213510 $Y=648685
X1192 57 369 5 4 365 AN2D1BWP7T $T=221640 703800 1 180 $X=218550 $Y=703565
X1193 388 369 5 4 382 AN2D1BWP7T $T=231720 743000 0 180 $X=228630 $Y=738790
X1194 310 314 5 4 340 AN2D1BWP7T $T=244040 641080 0 180 $X=240950 $Y=636870
X1195 364 82 5 4 404 AN2D1BWP7T $T=253560 625400 0 180 $X=250470 $Y=621190
X1196 388 261 5 4 444 AN2D1BWP7T $T=273720 735160 1 180 $X=270630 $Y=734925
X1197 456 82 5 4 461 AN2D1BWP7T $T=293320 648920 1 180 $X=290230 $Y=648685
X1198 473 82 5 4 459 AN2D1BWP7T $T=295560 641080 0 180 $X=292470 $Y=636870
X1199 456 479 5 4 405 AN2D1BWP7T $T=329720 711640 0 180 $X=326630 $Y=707430
X1200 568 82 5 4 496 AN2D1BWP7T $T=352680 719480 0 180 $X=349590 $Y=715270
X1201 121 119 5 4 118 AN2D1BWP7T $T=369480 609720 0 180 $X=366390 $Y=605510
X1202 121 480 5 4 618 AN2D1BWP7T $T=380120 601880 1 0 $X=379830 $Y=597670
X1203 516 482 5 4 603 AN2D1BWP7T $T=382360 648920 0 0 $X=382070 $Y=648685
X1204 144 119 5 4 654 AN2D1BWP7T $T=402520 664600 1 180 $X=399430 $Y=664365
X1205 179 119 5 4 662 AN2D1BWP7T $T=431640 601880 0 180 $X=428550 $Y=597670
X1206 338 331 406 4 5 411 XOR3D0BWP7T $T=244040 656760 1 0 $X=243750 $Y=652550
X1207 535 512 538 4 5 561 XOR3D0BWP7T $T=337560 601880 1 0 $X=337270 $Y=597670
X1208 304 317 315 4 5 393 XNR3D0BWP7T $T=225000 703800 1 0 $X=224710 $Y=699590
X1209 436 443 420 4 5 446 XNR3D0BWP7T $T=267000 633240 0 0 $X=266710 $Y=633005
X1210 99 484 100 4 5 476 XNR3D0BWP7T $T=307880 641080 1 180 $X=298070 $Y=640845
X1211 578 579 601 4 5 613 XNR3D0BWP7T $T=370600 609720 0 0 $X=370310 $Y=609485
X1212 304 315 5 363 311 4 IOA21D0BWP7T $T=215480 703800 0 0 $X=215190 $Y=703565
X1213 578 601 5 608 602 4 IOA21D0BWP7T $T=380120 648920 1 180 $X=376470 $Y=648685
X1214 478 5 108 467 4 510 109 OAI211D0BWP7T $T=328040 617560 1 0 $X=327750 $Y=613350
X1215 536 108 348 88 5 4 417 AO22D0BWP7T $T=336440 680280 1 180 $X=331670 $Y=680045
X1216 541 108 501 88 5 4 465 AO22D0BWP7T $T=338120 703800 1 180 $X=333350 $Y=703565
X1217 117 108 576 88 5 4 569 AO22D0BWP7T $T=360520 633240 0 180 $X=355750 $Y=629030
X1218 658 108 627 88 5 4 651 AO22D0BWP7T $T=402520 617560 0 180 $X=397750 $Y=613350
X1219 193 166 187 191 5 4 MAOI222D2BWP7T $T=444520 680280 1 180 $X=436950 $Y=680045
X1220 25 272 5 4 271 DFQD1BWP7T $T=180200 680280 0 0 $X=179910 $Y=680045
X1221 25 288 5 4 314 DFQD1BWP7T $T=225000 664600 1 180 $X=214070 $Y=664365
X1222 25 404 5 4 86 DFQD1BWP7T $T=265320 609720 0 180 $X=254390 $Y=605510
X1223 25 91 5 4 371 DFQD1BWP7T $T=276520 609720 0 180 $X=265590 $Y=605510
X1224 25 495 5 4 479 DFQD1BWP7T $T=312360 695960 0 180 $X=301430 $Y=691750
X1225 25 547 5 4 509 DFQD1BWP7T $T=343720 633240 1 180 $X=332790 $Y=633005
X1226 25 555 5 4 292 DFQD1BWP7T $T=347640 735160 1 180 $X=336710 $Y=734925
X1227 25 112 5 4 480 DFQD1BWP7T $T=352120 609720 1 180 $X=341190 $Y=609485
X1228 25 600 5 4 502 DFQD1BWP7T $T=377320 735160 1 180 $X=366390 $Y=734925
X1229 25 651 5 4 541 DFQD1BWP7T $T=402520 641080 1 180 $X=391590 $Y=640845
X1230 150 148 5 4 617 DFQD1BWP7T $T=419320 617560 1 180 $X=408390 $Y=617325
X1231 25 630 5 4 553 DFQD1BWP7T $T=419320 672440 1 180 $X=408390 $Y=672205
X1232 25 151 5 4 514 DFQD1BWP7T $T=422120 648920 0 180 $X=411190 $Y=644710
X1233 25 162 5 4 522 DFQD1BWP7T $T=429400 672440 0 180 $X=418470 $Y=668230
X1234 150 167 5 4 658 DFQD1BWP7T $T=430520 617560 1 180 $X=419590 $Y=617325
X1235 150 176 5 4 568 DFQD1BWP7T $T=433320 633240 0 180 $X=422390 $Y=629030
X1236 150 675 5 4 379 DFQD1BWP7T $T=443960 625400 0 180 $X=433030 $Y=621190
X1237 150 200 5 4 482 DFQD1BWP7T $T=443960 656760 0 180 $X=433030 $Y=652550
X1238 88 427 5 4 87 421 393 MOAI22D0BWP7T $T=262520 695960 0 180 $X=258310 $Y=691750
X1239 88 450 5 4 87 438 446 MOAI22D0BWP7T $T=276520 648920 1 180 $X=272310 $Y=648685
X1240 88 467 5 4 87 440 452 MOAI22D0BWP7T $T=295000 680280 0 180 $X=290790 $Y=676070
X1241 88 102 5 4 87 464 476 MOAI22D0BWP7T $T=302840 656760 1 180 $X=298630 $Y=656525
X1242 88 128 5 4 561 547 87 MOAI22D0BWP7T $T=374520 625400 1 180 $X=370310 $Y=625165
X1243 88 617 5 4 87 615 613 MOAI22D0BWP7T $T=382360 601880 1 180 $X=378150 $Y=601645
X1244 201 197 5 4 195 675 188 MOAI22D0BWP7T $T=441160 641080 1 180 $X=436950 $Y=640845
X1245 282 305 297 262 284 5 4 XNR4D0BWP7T $T=192520 648920 0 180 $X=179350 $Y=644710
X1246 297 357 54 367 339 5 4 XNR4D0BWP7T $T=211560 641080 1 0 $X=211270 $Y=636870
X1247 454 462 472 474 433 5 4 XNR4D0BWP7T $T=287720 719480 0 0 $X=287430 $Y=719245
X1248 472 551 542 523 457 5 4 XNR4D0BWP7T $T=345960 719480 0 180 $X=332790 $Y=715270
X1249 634 589 629 641 650 5 4 XNR4D0BWP7T $T=389080 680280 1 0 $X=388790 $Y=676070
X1250 636 643 634 642 657 5 4 XNR4D0BWP7T $T=389640 703800 0 0 $X=389350 $Y=703565
X1251 248 267 262 244 238 5 4 XOR4D0BWP7T $T=177400 664600 0 180 $X=164230 $Y=660390
X1252 325 274 339 341 346 5 4 XOR4D0BWP7T $T=198680 664600 1 0 $X=198390 $Y=660390
X1253 361 383 367 58 372 5 4 XOR4D0BWP7T $T=233400 625400 0 180 $X=220230 $Y=621190
X1254 414 412 457 373 432 5 4 XOR4D0BWP7T $T=297240 711640 0 180 $X=284070 $Y=707430
X1255 458 449 474 483 491 5 4 XOR4D0BWP7T $T=294440 735160 0 0 $X=294150 $Y=734925
X1256 526 530 523 503 439 5 4 XOR4D0BWP7T $T=337560 695960 1 180 $X=324390 $Y=695725
X1257 587 590 642 597 647 5 4 XOR4D0BWP7T $T=385160 664600 1 0 $X=384870 $Y=660390
X1258 621 649 641 624 633 5 4 XOR4D0BWP7T $T=401400 625400 1 180 $X=388230 $Y=625165
X1259 622 584 650 652 553 5 4 XOR4D0BWP7T $T=389640 688120 0 0 $X=389350 $Y=687885
X1260 64 5 4 60 CKND1BWP7T $T=228920 601880 1 180 $X=226950 $Y=601645
X1261 398 5 4 101 CKND1BWP7T $T=301720 609720 0 180 $X=299750 $Y=605510
X1262 591 5 4 528 CKND1BWP7T $T=421560 711640 0 180 $X=419590 $Y=707430
X1263 271 240 5 4 BUFFD1P5BWP7T $T=173480 711640 1 0 $X=173190 $Y=707430
X1264 502 261 5 4 BUFFD1P5BWP7T $T=314600 743000 0 180 $X=311510 $Y=738790
X1265 517 369 5 4 BUFFD1P5BWP7T $T=328040 719480 1 180 $X=324950 $Y=719245
X1266 275 4 232 428 5 NR2D0BWP7T $T=276520 711640 0 180 $X=273990 $Y=707430
X1267 37 320 4 296 5 35 319 AOI22D1BWP7T $T=192520 672440 1 180 $X=188310 $Y=672205
X1268 50 49 4 45 5 43 270 AOI22D1BWP7T $T=216600 680280 1 180 $X=212390 $Y=680045
X1269 37 353 4 283 5 35 286 AOI22D1BWP7T $T=221080 695960 1 180 $X=216870 $Y=695725
X1270 56 49 4 52 5 43 294 AOI22D1BWP7T $T=221640 680280 1 180 $X=217430 $Y=680045
X1271 37 374 4 371 5 35 266 AOI22D1BWP7T $T=222760 695960 0 180 $X=218550 $Y=691750
X1272 37 373 4 341 5 35 377 AOI22D1BWP7T $T=219960 688120 0 0 $X=219670 $Y=687885
X1273 37 256 4 46 5 35 378 AOI22D1BWP7T $T=229480 609720 1 180 $X=225270 $Y=609485
X1274 71 49 4 63 5 43 380 AOI22D1BWP7T $T=230040 680280 1 180 $X=225830 $Y=680045
X1275 77 49 4 75 5 43 381 AOI22D1BWP7T $T=249640 633240 1 180 $X=245430 $Y=633005
X1276 219 5 4 249 CKBD1BWP7T $T=162280 680280 0 0 $X=161990 $Y=680045
X1277 401 5 4 256 CKBD1BWP7T $T=246280 680280 0 0 $X=245990 $Y=680045
X1278 419 5 4 24 CKBD1BWP7T $T=258040 625400 1 180 $X=255510 $Y=625165
X1279 422 5 4 374 CKBD1BWP7T $T=259160 656760 0 0 $X=258870 $Y=656525
X1280 451 5 4 320 CKBD1BWP7T $T=282680 672440 1 0 $X=282390 $Y=668230
X1281 453 5 4 57 CKBD1BWP7T $T=286040 695960 1 0 $X=285750 $Y=691750
X1282 475 5 4 388 CKBD1BWP7T $T=296680 703800 0 0 $X=296390 $Y=703565
X1283 492 5 4 295 CKBD1BWP7T $T=305640 727320 1 0 $X=305350 $Y=723110
X1284 500 5 4 228 CKBD1BWP7T $T=313480 735160 0 180 $X=310950 $Y=730950
X1285 493 5 4 312 CKBD1BWP7T $T=326920 719480 1 0 $X=326630 $Y=715270
X1286 529 5 4 442 CKBD1BWP7T $T=334200 727320 1 180 $X=331670 $Y=727085
X1287 571 5 4 473 CKBD1BWP7T $T=354920 719480 0 180 $X=352390 $Y=715270
X1288 585 5 4 456 CKBD1BWP7T $T=368920 711640 1 180 $X=366390 $Y=711405
X1289 593 5 4 594 CKBD1BWP7T $T=368920 617560 0 0 $X=368630 $Y=617325
X1290 609 5 4 27 CKBD1BWP7T $T=376760 735160 1 0 $X=376470 $Y=730950
X1291 619 5 4 591 CKBD1BWP7T $T=381800 617560 0 0 $X=381510 $Y=617325
X1292 632 5 4 448 CKBD1BWP7T $T=387960 735160 0 0 $X=387670 $Y=734925
X1293 660 5 4 516 CKBD1BWP7T $T=413160 680280 1 180 $X=410630 $Y=680045
X1294 626 5 4 427 CKBD1BWP7T $T=415400 680280 1 180 $X=412870 $Y=680045
X1295 560 543 5 4 INVD1P5BWP7T $T=360520 664600 1 180 $X=357990 $Y=664365
X1296 564 30 5 4 INVD1P5BWP7T $T=414840 735160 1 180 $X=412310 $Y=734925
X1297 296 287 282 4 5 281 OA21D0BWP7T $T=182440 703800 0 180 $X=178790 $Y=699590
X1298 76 78 80 4 5 84 OA21D0BWP7T $T=249640 609720 1 0 $X=249350 $Y=605510
X1299 320 444 454 4 5 426 OA21D0BWP7T $T=285480 735160 1 0 $X=285190 $Y=730950
X1300 658 656 147 4 5 661 OA21D0BWP7T $T=413720 609720 0 0 $X=413430 $Y=609485
X1301 541 527 636 4 5 653 OA21D0BWP7T $T=421560 711640 1 0 $X=421270 $Y=707430
X1302 366 356 35 37 36 4 5 AOI22D0BWP7T $T=219400 656760 0 180 $X=215750 $Y=652550
X1303 370 368 35 37 362 4 5 AOI22D0BWP7T $T=221080 664600 0 180 $X=217430 $Y=660390
X1304 49 386 43 379 62 4 5 AOI22D0BWP7T $T=231160 672440 1 180 $X=227510 $Y=672205
X1305 49 385 43 70 68 4 5 AOI22D0BWP7T $T=233960 633240 1 180 $X=230310 $Y=633005
X1306 302 399 35 37 73 4 5 AOI22D0BWP7T $T=245720 609720 1 180 $X=242070 $Y=609485
X1307 49 415 43 83 81 4 5 AOI22D0BWP7T $T=255240 601880 0 180 $X=251590 $Y=597670
X1308 103 4 25 5 CKND10BWP7T $T=309560 648920 0 0 $X=309270 $Y=648685
X1309 5 4 ICV_76 $T=155000 688120 0 0 $X=154710 $Y=687885
X1310 5 4 ICV_76 $T=155000 695960 0 0 $X=154710 $Y=695725
X1311 5 4 ICV_76 $T=155000 703800 1 0 $X=154710 $Y=699590
X1312 5 4 ICV_76 $T=155000 735160 0 0 $X=154710 $Y=734925
X1313 5 4 ICV_76 $T=197000 688120 0 0 $X=196710 $Y=687885
X1314 5 4 ICV_76 $T=197000 695960 0 0 $X=196710 $Y=695725
X1315 5 4 ICV_76 $T=197000 719480 1 0 $X=196710 $Y=715270
X1316 5 4 ICV_76 $T=239000 648920 0 0 $X=238710 $Y=648685
X1317 5 4 ICV_76 $T=239000 688120 1 0 $X=238710 $Y=683910
X1318 5 4 ICV_76 $T=281000 609720 1 0 $X=280710 $Y=605510
X1319 5 4 ICV_76 $T=281000 617560 0 0 $X=280710 $Y=617325
X1320 5 4 ICV_76 $T=281000 633240 0 0 $X=280710 $Y=633005
X1321 5 4 ICV_76 $T=323000 609720 1 0 $X=322710 $Y=605510
X1322 5 4 ICV_76 $T=365000 617560 1 0 $X=364710 $Y=613350
X1323 5 4 ICV_76 $T=407000 601880 0 0 $X=406710 $Y=601645
X1324 5 4 ICV_76 $T=407000 609720 1 0 $X=406710 $Y=605510
X1325 5 4 ICV_76 $T=407000 617560 1 0 $X=406710 $Y=613350
X1326 5 4 ICV_76 $T=407000 664600 0 0 $X=406710 $Y=664365
X1327 5 4 ICV_41 $T=181880 648920 0 0 $X=181590 $Y=648685
X1328 5 4 ICV_41 $T=182440 711640 1 0 $X=182150 $Y=707430
X1329 5 4 ICV_41 $T=198120 617560 1 0 $X=197830 $Y=613350
X1330 5 4 ICV_41 $T=198120 641080 1 0 $X=197830 $Y=636870
X1331 5 4 ICV_41 $T=198120 680280 0 0 $X=197830 $Y=680045
X1332 5 4 ICV_41 $T=211560 601880 0 0 $X=211270 $Y=601645
X1333 5 4 ICV_41 $T=224440 641080 1 0 $X=224150 $Y=636870
X1334 5 4 ICV_41 $T=224440 719480 0 0 $X=224150 $Y=719245
X1335 5 4 ICV_41 $T=240120 617560 1 0 $X=239830 $Y=613350
X1336 5 4 ICV_41 $T=240120 617560 0 0 $X=239830 $Y=617325
X1337 5 4 ICV_41 $T=258040 735160 1 0 $X=257750 $Y=730950
X1338 5 4 ICV_41 $T=282120 703800 0 0 $X=281830 $Y=703565
X1339 5 4 ICV_41 $T=307880 641080 0 0 $X=307590 $Y=640845
X1340 5 4 ICV_41 $T=307880 719480 1 0 $X=307590 $Y=715270
X1341 5 4 ICV_41 $T=309000 680280 1 0 $X=308710 $Y=676070
X1342 5 4 ICV_41 $T=309560 703800 0 0 $X=309270 $Y=703565
X1343 5 4 ICV_41 $T=369480 609720 1 0 $X=369190 $Y=605510
X1344 5 4 ICV_41 $T=391880 688120 1 0 $X=391590 $Y=683910
X1345 5 4 ICV_41 $T=408120 688120 1 0 $X=407830 $Y=683910
X1346 5 4 ICV_41 $T=408120 688120 0 0 $X=407830 $Y=687885
X1347 5 4 ICV_41 $T=408120 703800 1 0 $X=407830 $Y=699590
X1348 5 4 ICV_41 $T=426040 617560 1 0 $X=425750 $Y=613350
X1349 5 4 ICV_41 $T=433880 648920 1 0 $X=433590 $Y=644710
X1350 5 4 ICV_41 $T=433880 672440 0 0 $X=433590 $Y=672205
X1351 5 4 ICV_37 $T=156120 601880 1 0 $X=155830 $Y=597670
X1352 5 4 ICV_37 $T=156120 648920 1 0 $X=155830 $Y=644710
X1353 5 4 ICV_37 $T=156120 648920 0 0 $X=155830 $Y=648685
X1354 5 4 ICV_37 $T=156120 672440 1 0 $X=155830 $Y=668230
X1355 5 4 ICV_37 $T=156120 727320 1 0 $X=155830 $Y=723110
X1356 5 4 ICV_37 $T=162840 735160 1 0 $X=162550 $Y=730950
X1357 5 4 ICV_37 $T=174600 672440 0 0 $X=174310 $Y=672205
X1358 5 4 ICV_37 $T=179640 601880 0 0 $X=179350 $Y=601645
X1359 5 4 ICV_37 $T=183000 672440 0 0 $X=182710 $Y=672205
X1360 5 4 ICV_37 $T=184680 703800 0 0 $X=184390 $Y=703565
X1361 5 4 ICV_37 $T=193640 617560 1 0 $X=193350 $Y=613350
X1362 5 4 ICV_37 $T=198120 680280 1 0 $X=197830 $Y=676070
X1363 5 4 ICV_37 $T=207080 609720 0 0 $X=206790 $Y=609485
X1364 5 4 ICV_37 $T=224440 672440 0 0 $X=224150 $Y=672205
X1365 5 4 ICV_37 $T=225000 664600 0 0 $X=224710 $Y=664365
X1366 5 4 ICV_37 $T=235640 672440 0 0 $X=235350 $Y=672205
X1367 5 4 ICV_37 $T=262520 625400 1 0 $X=262230 $Y=621190
X1368 5 4 ICV_37 $T=282120 656760 1 0 $X=281830 $Y=652550
X1369 5 4 ICV_37 $T=282120 735160 1 0 $X=281830 $Y=730950
X1370 5 4 ICV_37 $T=282120 735160 0 0 $X=281830 $Y=734925
X1371 5 4 ICV_37 $T=298920 680280 0 0 $X=298630 $Y=680045
X1372 5 4 ICV_37 $T=300040 719480 1 0 $X=299750 $Y=715270
X1373 5 4 ICV_37 $T=312920 625400 1 0 $X=312630 $Y=621190
X1374 5 4 ICV_37 $T=345960 719480 1 0 $X=345670 $Y=715270
X1375 5 4 ICV_37 $T=354920 641080 0 0 $X=354630 $Y=640845
X1376 5 4 ICV_37 $T=372280 601880 1 0 $X=371990 $Y=597670
X1377 5 4 ICV_37 $T=375080 601880 0 0 $X=374790 $Y=601645
X1378 5 4 ICV_37 $T=375080 648920 1 0 $X=374790 $Y=644710
X1379 5 4 ICV_37 $T=386280 719480 0 0 $X=385990 $Y=719245
X1380 5 4 ICV_37 $T=403640 617560 0 0 $X=403350 $Y=617325
X1381 5 4 ICV_37 $T=408120 648920 1 0 $X=407830 $Y=644710
X1382 5 4 ICV_37 $T=428280 672440 0 0 $X=427990 $Y=672205
X1383 5 4 ICV_37 $T=428280 735160 0 0 $X=427990 $Y=734925
X1384 5 4 ICV_37 $T=435000 664600 1 0 $X=434710 $Y=660390
X1385 5 4 ICV_37 $T=438920 609720 1 0 $X=438630 $Y=605510
X1386 5 4 ICV_37 $T=445640 641080 0 0 $X=445350 $Y=640845
X1387 5 4 ICV_37 $T=445640 703800 1 0 $X=445350 $Y=699590
X1388 5 4 ICV_60 $T=165080 633240 0 0 $X=164790 $Y=633005
X1389 5 4 ICV_60 $T=174040 703800 1 0 $X=173750 $Y=699590
X1390 5 4 ICV_60 $T=181320 719480 1 0 $X=181030 $Y=715270
X1391 5 4 ICV_60 $T=207080 735160 1 0 $X=206790 $Y=730950
X1392 5 4 ICV_60 $T=258040 688120 1 0 $X=257750 $Y=683910
X1393 5 4 ICV_60 $T=282120 664600 1 0 $X=281830 $Y=660390
X1394 5 4 ICV_60 $T=305080 656760 1 0 $X=304790 $Y=652550
X1395 5 4 ICV_60 $T=309000 672440 0 0 $X=308710 $Y=672205
X1396 5 4 ICV_60 $T=309000 688120 1 0 $X=308710 $Y=683910
X1397 5 4 ICV_60 $T=351000 617560 1 0 $X=350710 $Y=613350
X1398 5 4 ICV_60 $T=351000 633240 1 0 $X=350710 $Y=629030
X1399 5 4 ICV_60 $T=368920 641080 0 0 $X=368630 $Y=640845
X1400 5 4 ICV_60 $T=393000 617560 1 0 $X=392710 $Y=613350
X1401 5 4 ICV_60 $T=423800 711640 0 0 $X=423510 $Y=711405
X1402 5 4 ICV_60 $T=443960 625400 1 0 $X=443670 $Y=621190
X1403 5 4 ICV_60 $T=443960 633240 0 0 $X=443670 $Y=633005
X1404 5 4 ICV_60 $T=443960 648920 0 0 $X=443670 $Y=648685
X1405 5 4 ICV_60 $T=443960 656760 1 0 $X=443670 $Y=652550
X1406 5 4 ICV_60 $T=443960 695960 1 0 $X=443670 $Y=691750
X1407 5 4 ICV_60 $T=443960 695960 0 0 $X=443670 $Y=695725
X1408 5 4 ICV_60 $T=443960 703800 0 0 $X=443670 $Y=703565
X1409 5 4 ICV_60 $T=443960 719480 1 0 $X=443670 $Y=715270
X1410 5 4 ICV_60 $T=443960 743000 1 0 $X=443670 $Y=738790
X1411 5 4 ICV_43 $T=176280 719480 1 0 $X=175990 $Y=715270
X1412 5 4 ICV_43 $T=177400 735160 0 0 $X=177110 $Y=734925
X1413 5 4 ICV_43 $T=217720 625400 1 0 $X=217430 $Y=621190
X1414 5 4 ICV_43 $T=249080 601880 1 0 $X=248790 $Y=597670
X1415 5 4 ICV_43 $T=249080 727320 1 0 $X=248790 $Y=723110
X1416 5 4 ICV_43 $T=253000 625400 0 0 $X=252710 $Y=625165
X1417 5 4 ICV_43 $T=258040 648920 0 0 $X=257750 $Y=648685
X1418 5 4 ICV_43 $T=266440 735160 0 0 $X=266150 $Y=734925
X1419 5 4 ICV_43 $T=269800 648920 0 0 $X=269510 $Y=648685
X1420 5 4 ICV_43 $T=282120 641080 0 0 $X=281830 $Y=640845
X1421 5 4 ICV_43 $T=285480 680280 0 0 $X=285190 $Y=680045
X1422 5 4 ICV_43 $T=291080 601880 1 0 $X=290790 $Y=597670
X1423 5 4 ICV_43 $T=295560 641080 0 0 $X=295270 $Y=640845
X1424 5 4 ICV_43 $T=298920 695960 1 0 $X=298630 $Y=691750
X1425 5 4 ICV_43 $T=309000 743000 1 0 $X=308710 $Y=738790
X1426 5 4 ICV_43 $T=324120 641080 0 0 $X=323830 $Y=640845
X1427 5 4 ICV_43 $T=324120 664600 1 0 $X=323830 $Y=660390
X1428 5 4 ICV_43 $T=324120 719480 1 0 $X=323830 $Y=715270
X1429 5 4 ICV_43 $T=327480 664600 0 0 $X=327190 $Y=664365
X1430 5 4 ICV_43 $T=329720 656760 1 0 $X=329430 $Y=652550
X1431 5 4 ICV_43 $T=342040 680280 1 0 $X=341750 $Y=676070
X1432 5 4 ICV_43 $T=366120 672440 0 0 $X=365830 $Y=672205
X1433 5 4 ICV_43 $T=370600 648920 0 0 $X=370310 $Y=648685
X1434 5 4 ICV_43 $T=375080 727320 1 0 $X=374790 $Y=723110
X1435 5 4 ICV_43 $T=408120 680280 0 0 $X=407830 $Y=680045
X1436 5 4 ICV_43 $T=419320 680280 0 0 $X=419030 $Y=680045
X1437 5 4 ICV_43 $T=446200 680280 1 0 $X=445910 $Y=676070
X1438 5 4 ICV_43 $T=446200 688120 0 0 $X=445910 $Y=687885
X1439 5 4 ICV_52 $T=156120 641080 1 0 $X=155830 $Y=636870
X1440 5 4 ICV_52 $T=156120 641080 0 0 $X=155830 $Y=640845
X1441 5 4 ICV_52 $T=216040 688120 0 0 $X=215750 $Y=687885
X1442 5 4 ICV_52 $T=240120 648920 1 0 $X=239830 $Y=644710
X1443 5 4 ICV_52 $T=240120 656760 1 0 $X=239830 $Y=652550
X1444 5 4 ICV_52 $T=277080 680280 0 0 $X=276790 $Y=680045
X1445 5 4 ICV_52 $T=282120 695960 1 0 $X=281830 $Y=691750
X1446 5 4 ICV_52 $T=290520 735160 0 0 $X=290230 $Y=734925
X1447 5 4 ICV_52 $T=301720 609720 1 0 $X=301430 $Y=605510
X1448 5 4 ICV_52 $T=329160 719480 1 0 $X=328870 $Y=715270
X1449 5 4 ICV_52 $T=361080 609720 0 0 $X=360790 $Y=609485
X1450 5 4 ICV_52 $T=375080 688120 1 0 $X=374790 $Y=683910
X1451 5 4 ICV_52 $T=381240 633240 0 0 $X=380950 $Y=633005
X1452 5 4 ICV_52 $T=395800 656760 1 0 $X=395510 $Y=652550
X1453 5 4 ICV_52 $T=395800 664600 0 0 $X=395510 $Y=664365
X1454 5 4 ICV_52 $T=403080 719480 1 0 $X=402790 $Y=715270
X1455 5 4 ICV_52 $T=408120 601880 1 0 $X=407830 $Y=597670
X1456 5 4 ICV_52 $T=421560 695960 0 0 $X=421270 $Y=695725
X1457 5 4 ICV_52 $T=424920 601880 1 0 $X=424630 $Y=597670
X1458 5 4 ICV_52 $T=445080 656760 0 0 $X=444790 $Y=656525
X1459 5 4 ICV_54 $T=213240 695960 1 0 $X=212950 $Y=691750
X1460 5 4 ICV_54 $T=216040 719480 1 0 $X=215750 $Y=715270
X1461 5 4 ICV_54 $T=219960 609720 0 0 $X=219670 $Y=609485
X1462 5 4 ICV_54 $T=233400 625400 1 0 $X=233110 $Y=621190
X1463 5 4 ICV_54 $T=233400 735160 0 0 $X=233110 $Y=734925
X1464 5 4 ICV_54 $T=240120 633240 0 0 $X=239830 $Y=633005
X1465 5 4 ICV_54 $T=254680 648920 1 0 $X=254390 $Y=644710
X1466 5 4 ICV_54 $T=282120 719480 0 0 $X=281830 $Y=719245
X1467 5 4 ICV_54 $T=300040 633240 0 0 $X=299750 $Y=633005
X1468 5 4 ICV_54 $T=317400 695960 0 0 $X=317110 $Y=695725
X1469 5 4 ICV_54 $T=324120 609720 0 0 $X=323830 $Y=609485
X1470 5 4 ICV_54 $T=359400 680280 1 0 $X=359110 $Y=676070
X1471 5 4 ICV_54 $T=368920 711640 0 0 $X=368630 $Y=711405
X1472 5 4 ICV_54 $T=391320 601880 0 0 $X=391030 $Y=601645
X1473 5 4 ICV_54 $T=408120 609720 0 0 $X=407830 $Y=609485
X1474 5 4 ICV_54 $T=413720 711640 0 0 $X=413430 $Y=711405
X1475 5 4 ICV_54 $T=427160 688120 1 0 $X=426870 $Y=683910
X1476 5 4 ICV_54 $T=429400 672440 1 0 $X=429110 $Y=668230
X1477 5 4 ICV_38 $T=192520 703800 0 0 $X=192230 $Y=703565
X1478 5 4 ICV_38 $T=234520 719480 1 0 $X=234230 $Y=715270
X1479 5 4 ICV_38 $T=276520 648920 0 0 $X=276230 $Y=648685
X1480 5 4 ICV_38 $T=276520 664600 0 0 $X=276230 $Y=664365
X1481 5 4 ICV_38 $T=276520 711640 1 0 $X=276230 $Y=707430
X1482 5 4 ICV_38 $T=276520 719480 0 0 $X=276230 $Y=719245
X1483 5 4 ICV_38 $T=318520 633240 0 0 $X=318230 $Y=633005
X1484 5 4 ICV_38 $T=318520 719480 0 0 $X=318230 $Y=719245
X1485 5 4 ICV_38 $T=318520 727320 1 0 $X=318230 $Y=723110
X1486 5 4 ICV_38 $T=360520 633240 1 0 $X=360230 $Y=629030
X1487 5 4 ICV_38 $T=360520 695960 1 0 $X=360230 $Y=691750
X1488 5 4 ICV_38 $T=402520 641080 0 0 $X=402230 $Y=640845
X1489 5 4 ICV_38 $T=402520 656760 0 0 $X=402230 $Y=656525
X1490 5 4 ICV_38 $T=402520 688120 0 0 $X=402230 $Y=687885
X1491 5 4 ICV_38 $T=402520 703800 0 0 $X=402230 $Y=703565
X1492 5 4 ICV_38 $T=402520 719480 0 0 $X=402230 $Y=719245
X1493 5 4 ICV_45 $T=162280 601880 1 0 $X=161990 $Y=597670
X1494 5 4 ICV_45 $T=162280 641080 0 0 $X=161990 $Y=640845
X1495 5 4 ICV_45 $T=162840 680280 1 0 $X=162550 $Y=676070
X1496 5 4 ICV_45 $T=198120 609720 1 0 $X=197830 $Y=605510
X1497 5 4 ICV_45 $T=198120 703800 1 0 $X=197830 $Y=699590
X1498 5 4 ICV_45 $T=282120 672440 0 0 $X=281830 $Y=672205
X1499 5 4 ICV_45 $T=282120 688120 1 0 $X=281830 $Y=683910
X1500 5 4 ICV_45 $T=282120 743000 1 0 $X=281830 $Y=738790
X1501 5 4 ICV_45 $T=293320 601880 0 0 $X=293030 $Y=601645
X1502 5 4 ICV_45 $T=293320 617560 1 0 $X=293030 $Y=613350
X1503 5 4 ICV_45 $T=324120 633240 1 0 $X=323830 $Y=629030
X1504 5 4 ICV_45 $T=337560 625400 0 0 $X=337270 $Y=625165
X1505 5 4 ICV_45 $T=337560 695960 0 0 $X=337270 $Y=695725
X1506 5 4 ICV_45 $T=368920 656760 1 0 $X=368630 $Y=652550
X1507 5 4 ICV_45 $T=380120 609720 0 0 $X=379830 $Y=609485
X1508 5 4 ICV_45 $T=408120 625400 0 0 $X=407830 $Y=625165
X1509 145 5 4 659 BUFFD1BWP7T $T=411480 641080 1 180 $X=408950 $Y=640845
X1510 617 639 5 4 645 137 IAO21D0BWP7T $T=391880 601880 1 0 $X=391590 $Y=597670
X1511 522 560 509 4 5 525 AN3D1BWP7T $T=353800 680280 1 0 $X=353510 $Y=676070
X1512 522 595 536 4 5 586 AN3D1BWP7T $T=386840 711640 1 180 $X=383190 $Y=711405
X1513 138 140 617 4 5 645 AN3D1BWP7T $T=396920 601880 0 0 $X=396630 $Y=601645
X1514 522 594 427 4 5 644 AN3D1BWP7T $T=410360 711640 0 0 $X=410070 $Y=711405
X1515 378 61 59 5 4 ND2D2BWP7T $T=225560 609720 1 0 $X=225270 $Y=605510
X1516 381 5 377 66 4 CKND2D2BWP7T $T=228360 648920 1 0 $X=228070 $Y=644710
X1517 5 4 ICV_69 $T=155000 601880 0 0 $X=154710 $Y=601645
X1518 5 4 ICV_69 $T=155000 672440 0 0 $X=154710 $Y=672205
X1519 5 4 ICV_69 $T=155000 688120 1 0 $X=154710 $Y=683910
X1520 5 4 ICV_69 $T=155000 711640 1 0 $X=154710 $Y=707430
X1521 5 4 ICV_69 $T=155000 711640 0 0 $X=154710 $Y=711405
X1522 5 4 ICV_69 $T=197000 601880 1 0 $X=196710 $Y=597670
X1523 5 4 ICV_69 $T=197000 625400 0 0 $X=196710 $Y=625165
X1524 5 4 ICV_69 $T=197000 648920 0 0 $X=196710 $Y=648685
X1525 5 4 ICV_69 $T=197000 735160 1 0 $X=196710 $Y=730950
X1526 5 4 ICV_69 $T=239000 601880 1 0 $X=238710 $Y=597670
X1527 5 4 ICV_69 $T=239000 664600 0 0 $X=238710 $Y=664365
X1528 5 4 ICV_69 $T=239000 695960 0 0 $X=238710 $Y=695725
X1529 5 4 ICV_69 $T=281000 601880 1 0 $X=280710 $Y=597670
X1530 5 4 ICV_69 $T=281000 609720 0 0 $X=280710 $Y=609485
X1531 5 4 ICV_69 $T=281000 625400 1 0 $X=280710 $Y=621190
X1532 5 4 ICV_69 $T=281000 641080 1 0 $X=280710 $Y=636870
X1533 5 4 ICV_69 $T=281000 656760 0 0 $X=280710 $Y=656525
X1534 5 4 ICV_69 $T=323000 625400 1 0 $X=322710 $Y=621190
X1535 5 4 ICV_69 $T=323000 695960 1 0 $X=322710 $Y=691750
X1536 5 4 ICV_69 $T=323000 703800 0 0 $X=322710 $Y=703565
X1537 5 4 ICV_69 $T=365000 648920 1 0 $X=364710 $Y=644710
X1538 5 4 ICV_69 $T=407000 641080 1 0 $X=406710 $Y=636870
X1539 88 485 5 434 397 87 4 MOAI22D1BWP7T $T=318520 672440 1 180 $X=313750 $Y=672205
X1540 88 553 5 87 470 542 4 MOAI22D1BWP7T $T=345400 680280 1 180 $X=340630 $Y=680045
X1541 88 136 5 87 630 629 4 MOAI22D1BWP7T $T=391320 648920 1 180 $X=386550 $Y=648685
X1542 509 582 4 525 531 5 IAO21D1BWP7T $T=366680 664600 1 0 $X=366390 $Y=660390
X1543 536 596 4 586 532 5 IAO21D1BWP7T $T=369480 703800 1 0 $X=369190 $Y=699590
X1544 427 607 4 644 605 5 IAO21D1BWP7T $T=403080 735160 0 180 $X=398870 $Y=730950
X1545 88 509 396 87 4 411 5 IOA22D2BWP7T $T=320200 688120 0 180 $X=313750 $Y=683910
X1546 88 113 504 87 4 534 5 IOA22D2BWP7T $T=356600 601880 0 180 $X=350150 $Y=597670
X1547 13 88 37 5 4 INR2XD4BWP7T $T=318520 609720 0 180 $X=305350 $Y=605510
X1548 371 5 42 314 4 398 ND3D1BWP7T $T=240680 625400 0 0 $X=240390 $Y=625165
X1549 374 5 479 369 4 418 ND3D1BWP7T $T=329720 680280 1 180 $X=326070 $Y=680045
X1550 50 5 161 202 4 194 ND3D1BWP7T $T=438920 688120 1 0 $X=438630 $Y=683910
X1551 5 4 ICV_75 $T=165080 711640 1 0 $X=164790 $Y=707430
X1552 5 4 ICV_75 $T=188600 727320 1 0 $X=188310 $Y=723110
X1553 5 4 ICV_75 $T=230600 664600 0 0 $X=230310 $Y=664365
X1554 5 4 ICV_75 $T=272600 609720 0 0 $X=272310 $Y=609485
X1555 5 4 ICV_75 $T=282120 648920 0 0 $X=281830 $Y=648685
X1556 5 4 ICV_75 $T=307320 664600 1 0 $X=307030 $Y=660390
X1557 5 4 ICV_75 $T=314600 672440 1 0 $X=314310 $Y=668230
X1558 5 4 ICV_75 $T=314600 743000 1 0 $X=314310 $Y=738790
X1559 5 4 ICV_75 $T=333080 625400 1 0 $X=332790 $Y=621190
X1560 5 4 ICV_75 $T=356600 601880 1 0 $X=356310 $Y=597670
X1561 5 4 ICV_75 $T=356600 625400 1 0 $X=356310 $Y=621190
X1562 5 4 ICV_75 $T=381240 703800 0 0 $X=380950 $Y=703565
X1563 5 4 ICV_75 $T=398600 648920 1 0 $X=398310 $Y=644710
X1564 5 4 ICV_75 $T=398600 648920 0 0 $X=398310 $Y=648685
X1565 5 4 ICV_75 $T=440600 664600 1 0 $X=440310 $Y=660390
X1566 5 4 ICV_75 $T=440600 727320 1 0 $X=440310 $Y=723110
X1567 5 4 ICV_74 $T=167880 719480 1 0 $X=167590 $Y=715270
X1568 5 4 ICV_74 $T=190840 680280 0 0 $X=190550 $Y=680045
X1569 5 4 ICV_74 $T=211560 664600 1 0 $X=211270 $Y=660390
X1570 5 4 ICV_74 $T=232840 617560 1 0 $X=232550 $Y=613350
X1571 5 4 ICV_74 $T=240120 680280 0 0 $X=239830 $Y=680045
X1572 5 4 ICV_74 $T=274840 641080 1 0 $X=274550 $Y=636870
X1573 5 4 ICV_74 $T=293320 633240 1 0 $X=293030 $Y=629030
X1574 5 4 ICV_74 $T=295560 672440 1 0 $X=295270 $Y=668230
X1575 5 4 ICV_74 $T=316840 648920 0 0 $X=316550 $Y=648685
X1576 5 4 ICV_74 $T=316840 695960 1 0 $X=316550 $Y=691750
X1577 5 4 ICV_74 $T=332520 641080 0 0 $X=332230 $Y=640845
X1578 5 4 ICV_74 $T=358840 648920 0 0 $X=358550 $Y=648685
X1579 5 4 ICV_74 $T=358840 703800 0 0 $X=358550 $Y=703565
X1580 5 4 ICV_74 $T=400840 735160 0 0 $X=400550 $Y=734925
X1581 5 4 ICV_74 $T=426040 601880 0 0 $X=425750 $Y=601645
X1582 5 4 ICV_74 $T=442840 711640 1 0 $X=442550 $Y=707430
X1583 36 300 4 33 34 5 OAI21D1BWP7T $T=189720 609720 0 180 $X=186070 $Y=605510
X1584 351 371 4 398 74 5 OAI21D1BWP7T $T=242920 601880 0 0 $X=242630 $Y=601645
X1585 485 487 4 489 494 5 OAI21D1BWP7T $T=303400 656760 0 0 $X=303110 $Y=656525
X1586 70 665 4 664 156 5 OAI21D1BWP7T $T=425480 680280 1 180 $X=421830 $Y=680045
.ENDS
***************************************
.SUBCKT ICV_33
** N=4 EP=0 IP=12 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_73 2 3 4 5 6 7 8 13 14
** N=18 EP=9 IP=128 FDC=410
*.SEEDPROM
X38 4 6 5 5 2 7 13 8 7 17 7 5 PDDW0208CDG $T=210000 900000 0 180 $X=129400 $Y=780000
X39 4 6 5 5 3 7 14 8 7 18 7 5 PDDW0208CDG $T=290030 900000 0 180 $X=209430 $Y=780000
X40 4 5 5 5 PVDD2CDG $T=370065 900000 0 180 $X=289465 $Y=780000
X41 4 5 PVSS3CDG $T=450100 900000 0 180 $X=369500 $Y=780000
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5 6 7
** N=9 EP=7 IP=13 FDC=145
*.SEEDPROM
X0 1 2 3 3 7 5 4 6 5 9 5 3 PDDW0208CDG $T=0 0 0 0 $X=-600 $Y=0
.ENDS
***************************************
.SUBCKT ICV_25 1 2 3 4 5 6 7
** N=9 EP=7 IP=13 FDC=145
*.SEEDPROM
X0 1 2 3 3 7 4 5 6 4 9 4 3 PDDW0208CDG $T=0 0 0 0 $X=-600 $Y=0
.ENDS
***************************************
.SUBCKT ICV_23 1 3
** N=5 EP=2 IP=6 FDC=60
*.SEEDPROM
X0 1 3 3 3 PVDD2CDG $T=0 0 0 0 $X=-600 $Y=0
.ENDS
***************************************
.SUBCKT HBK183_PREDRV_GR_VDD1DYN_S
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT HBK183_NMOS_W26_L03_DYN_S
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_PREDRV_VDD1CDG_DYN_S 2 3 4 5
** N=5 EP=4 IP=60 FDC=26
*.SEEDPROM
M0 2 4 3 5 N L=3e-07 W=2.6e-05 $X=5440 $Y=5210 $D=0
M1 3 4 2 5 N L=3e-07 W=2.6e-05 $X=9400 $Y=5210 $D=0
M2 2 4 3 5 N L=3e-07 W=2.6e-05 $X=10920 $Y=5210 $D=0
M3 3 4 2 5 N L=3e-07 W=2.6e-05 $X=14880 $Y=5210 $D=0
M4 2 4 3 5 N L=3e-07 W=2.6e-05 $X=16400 $Y=5210 $D=0
M5 3 4 2 5 N L=3e-07 W=2.6e-05 $X=20360 $Y=5210 $D=0
M6 2 4 3 5 N L=3e-07 W=2.6e-05 $X=21880 $Y=5210 $D=0
M7 3 4 2 5 N L=3e-07 W=2.6e-05 $X=25840 $Y=5210 $D=0
M8 2 4 3 5 N L=3e-07 W=2.6e-05 $X=27360 $Y=5210 $D=0
M9 3 4 2 5 N L=3e-07 W=2.6e-05 $X=31320 $Y=5210 $D=0
M10 2 4 3 5 N L=3e-07 W=2.6e-05 $X=32840 $Y=5210 $D=0
M11 3 4 2 5 N L=3e-07 W=2.6e-05 $X=36800 $Y=5210 $D=0
M12 2 4 3 5 N L=3e-07 W=2.6e-05 $X=38320 $Y=5210 $D=0
M13 3 4 2 5 N L=3e-07 W=2.6e-05 $X=42280 $Y=5210 $D=0
M14 2 4 3 5 N L=3e-07 W=2.6e-05 $X=43800 $Y=5210 $D=0
M15 3 4 2 5 N L=3e-07 W=2.6e-05 $X=47760 $Y=5210 $D=0
M16 2 4 3 5 N L=3e-07 W=2.6e-05 $X=49280 $Y=5210 $D=0
M17 3 4 2 5 N L=3e-07 W=2.6e-05 $X=53240 $Y=5210 $D=0
M18 2 4 3 5 N L=3e-07 W=2.6e-05 $X=54760 $Y=5210 $D=0
M19 3 4 2 5 N L=3e-07 W=2.6e-05 $X=58720 $Y=5210 $D=0
M20 2 4 3 5 N L=3e-07 W=2.6e-05 $X=60240 $Y=5210 $D=0
M21 3 4 2 5 N L=3e-07 W=2.6e-05 $X=64200 $Y=5210 $D=0
M22 2 4 3 5 N L=3e-07 W=2.6e-05 $X=65720 $Y=5210 $D=0
M23 3 4 2 5 N L=3e-07 W=2.6e-05 $X=69680 $Y=5210 $D=0
M24 2 4 3 5 N L=3e-07 W=2.6e-05 $X=71200 $Y=5210 $D=0
M25 3 4 2 5 N L=3e-07 W=2.6e-05 $X=75160 $Y=5210 $D=0
.ENDS
***************************************
.SUBCKT HBK183_NMOS_W15_L6D3_DYN
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_14
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_PDIODE_BASE_S
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT HBK183_RES_03_DYN
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT PVDD1CDG VDDPST VDD VSSPST VSS 6
** N=8 EP=5 IP=38 FDC=55
*.SEEDPROM
M0 VSSPST 8 VSSPST 6 ND L=4.18e-06 W=1.5e-05 $X=5030 $Y=5590 $D=1
M1 7 8 VSSPST 6 ND L=2e-06 W=5e-06 $X=5045 $Y=25430 $D=1
M2 VSSPST 8 VSSPST 6 ND L=4.18e-06 W=1.5e-05 $X=10510 $Y=5590 $D=1
M3 VSSPST 8 VSSPST 6 ND L=4.18e-06 W=1.5e-05 $X=15990 $Y=5590 $D=1
M4 VSSPST 8 VSSPST 6 ND L=4.18e-06 W=1.5e-05 $X=21470 $Y=5590 $D=1
M5 VSSPST 8 VSSPST 6 ND L=4.18e-06 W=1.5e-05 $X=26950 $Y=5590 $D=1
M6 VSSPST 8 VSSPST 6 ND L=4.18e-06 W=1.5e-05 $X=32430 $Y=5590 $D=1
M7 VSSPST 8 VSSPST 6 ND L=4.18e-06 W=1.5e-05 $X=37910 $Y=5590 $D=1
M8 VSSPST 8 VSSPST 6 ND L=4.18e-06 W=1.5e-05 $X=43390 $Y=5590 $D=1
M9 VSSPST 8 VSSPST 6 ND L=4.18e-06 W=1.5e-05 $X=48870 $Y=5590 $D=1
M10 VSSPST 8 VSSPST 6 ND L=4.18e-06 W=1.5e-05 $X=54350 $Y=5590 $D=1
M11 VSSPST 8 VSSPST 6 ND L=4.18e-06 W=1.5e-05 $X=59830 $Y=5590 $D=1
M12 VSSPST 8 VSSPST 6 ND L=4.18e-06 W=1.5e-05 $X=65310 $Y=5590 $D=1
M13 VSSPST 8 VSSPST 6 ND L=4.18e-06 W=1.5e-05 $X=70790 $Y=5590 $D=1
D14 VDD VDDPST D1 AREA=5.48392e-11 PJ=4.90684e-05 $X=5900 $Y=51960 $D=29
D15 VDD VDDPST D1 AREA=5.48392e-11 PJ=4.90684e-05 $X=11380 $Y=51960 $D=29
D16 VDD VDDPST D1 AREA=5.48392e-11 PJ=4.90684e-05 $X=16860 $Y=51960 $D=29
D17 VDD VDDPST D1 AREA=5.48392e-11 PJ=4.90684e-05 $X=22340 $Y=51960 $D=29
D18 VDD VDDPST D1 AREA=5.48392e-11 PJ=4.90684e-05 $X=27820 $Y=51960 $D=29
D19 VDD VDDPST D1 AREA=5.48392e-11 PJ=4.90684e-05 $X=33300 $Y=51960 $D=29
D20 VDD VDDPST D1 AREA=5.48392e-11 PJ=4.90684e-05 $X=38780 $Y=51960 $D=29
D21 VDD VDDPST D1 AREA=5.48392e-11 PJ=4.90684e-05 $X=44260 $Y=51960 $D=29
D22 VDD VDDPST D1 AREA=5.48392e-11 PJ=4.90684e-05 $X=49740 $Y=51960 $D=29
D23 VDD VDDPST D1 AREA=5.48392e-11 PJ=4.90684e-05 $X=55220 $Y=51960 $D=29
D24 VDD VDDPST D1 AREA=5.48392e-11 PJ=4.90684e-05 $X=60700 $Y=51960 $D=29
D25 VDD VDDPST D1 AREA=5.48392e-11 PJ=4.90684e-05 $X=66180 $Y=51960 $D=29
D26 VDD VDDPST D1 AREA=5.48392e-11 PJ=4.90684e-05 $X=71660 $Y=51960 $D=29
R27 8 VDD 1.0592e+06 $[PR] $X=9870 $Y=23910 $D=52
D28 6 VDDPST pnwdio_5_iso AREA=2.06895e-09 pj=0.0002054 $X=2410 $Y=49040 $D=112
X30 VDD VSS 7 6 HBK183_PREDRV_VDD1CDG_DYN_S $T=-450 80560 0 0 $X=-600 $Y=80410
.ENDS
***************************************
.SUBCKT ICV_18 1 2 3
** N=5 EP=3 IP=6 FDC=55
*.SEEDPROM
X0 1 2 3 3 3 PVDD1CDG $T=0 0 0 0 $X=-600 $Y=0
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3 4 5 6 7
** N=9 EP=7 IP=13 FDC=145
*.SEEDPROM
X0 1 2 3 3 7 5 4 6 5 9 5 3 PDDW0208CDG $T=0 0 0 0 $X=-600 $Y=0
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3 4 5 6 7
** N=9 EP=7 IP=13 FDC=145
*.SEEDPROM
X0 1 2 3 3 7 4 5 6 4 9 4 3 PDDW0208CDG $T=0 0 0 0 $X=-600 $Y=0
.ENDS
***************************************
.SUBCKT ICV_68 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=30
*.SEEDPROM
X0 1 2 DCAP8BWP7T $T=0 0 1 180 $X=-4770 $Y=-235
X1 3 4 1 2 5 DFQD0BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_35
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT INR2XD2BWP7T A1 B1 ZN VSS VDD
** N=10 EP=5 IP=0 FDC=14
*.SEEDPROM
M0 VSS A1 6 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 ZN 6 VSS VSS N L=1.8e-07 W=1e-06 $X=1470 $Y=345 $D=0
M2 VSS B1 ZN VSS N L=1.8e-07 W=1e-06 $X=2485 $Y=345 $D=0
M3 ZN B1 VSS VSS N L=1.8e-07 W=1e-06 $X=4400 $Y=345 $D=0
M4 VSS 6 ZN VSS N L=1.8e-07 W=1e-06 $X=5360 $Y=345 $D=0
M5 VDD A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M6 7 6 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1470 $Y=2205 $D=16
M7 ZN B1 7 VDD P L=1.8e-07 W=1.37e-06 $X=1910 $Y=2205 $D=16
M8 8 B1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2630 $Y=2205 $D=16
M9 VDD 6 8 VDD P L=1.8e-07 W=1.37e-06 $X=3060 $Y=2205 $D=16
M10 9 6 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3780 $Y=2205 $D=16
M11 ZN B1 9 VDD P L=1.8e-07 W=1.37e-06 $X=4210 $Y=2205 $D=16
M12 10 B1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4930 $Y=2205 $D=16
M13 VDD 6 10 VDD P L=1.8e-07 W=1.37e-06 $X=5360 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_70 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109
** N=352 EP=108 IP=3317 FDC=8130
*.SEEDPROM
M0 352 50 43 3 N L=1.8e-07 W=1e-06 $X=552715 $Y=233745 $D=0
M1 3 52 352 3 N L=1.8e-07 W=6.85e-07 $X=553440 $Y=233745 $D=0
M2 3 263 263 3 N L=1.8e-07 W=1e-06 $X=631200 $Y=161495 $D=0
M3 43 50 4 4 P L=1.8e-07 W=1.37e-06 $X=552715 $Y=235605 $D=16
M4 4 52 43 4 P L=1.8e-07 W=1.37e-06 $X=553440 $Y=235605 $D=16
M5 79 263 4 4 P L=1.8e-07 W=1.37e-06 $X=631200 $Y=159265 $D=16
X150 4 3 DCAPBWP7T $T=450120 209880 0 0 $X=449830 $Y=209645
X151 4 3 DCAPBWP7T $T=450120 233400 1 0 $X=449830 $Y=229190
X152 4 3 DCAPBWP7T $T=456840 155000 0 0 $X=456550 $Y=154765
X153 4 3 DCAPBWP7T $T=463560 202040 1 0 $X=463270 $Y=197830
X154 4 3 DCAPBWP7T $T=473640 178520 1 0 $X=473350 $Y=174310
X155 4 3 DCAPBWP7T $T=480920 241240 1 0 $X=480630 $Y=237030
X156 4 3 DCAPBWP7T $T=489320 186360 1 0 $X=489030 $Y=182150
X157 4 3 DCAPBWP7T $T=492120 194200 0 0 $X=491830 $Y=193965
X158 4 3 DCAPBWP7T $T=496600 202040 1 0 $X=496310 $Y=197830
X159 4 3 DCAPBWP7T $T=503880 162840 1 0 $X=503590 $Y=158630
X160 4 3 DCAPBWP7T $T=506120 209880 1 0 $X=505830 $Y=205670
X161 4 3 DCAPBWP7T $T=507800 225560 1 0 $X=507510 $Y=221350
X162 4 3 DCAPBWP7T $T=518440 225560 1 0 $X=518150 $Y=221350
X163 4 3 DCAPBWP7T $T=521240 178520 1 0 $X=520950 $Y=174310
X164 4 3 DCAPBWP7T $T=531320 170680 1 0 $X=531030 $Y=166470
X165 4 3 DCAPBWP7T $T=531320 178520 1 0 $X=531030 $Y=174310
X166 4 3 DCAPBWP7T $T=531320 194200 1 0 $X=531030 $Y=189990
X167 4 3 DCAPBWP7T $T=531320 194200 0 0 $X=531030 $Y=193965
X168 4 3 DCAPBWP7T $T=531320 233400 1 0 $X=531030 $Y=229190
X169 4 3 DCAPBWP7T $T=531320 241240 1 0 $X=531030 $Y=237030
X170 4 3 DCAPBWP7T $T=556520 217720 0 0 $X=556230 $Y=217485
X171 4 3 DCAPBWP7T $T=562680 178520 1 0 $X=562390 $Y=174310
X172 4 3 DCAPBWP7T $T=563800 202040 0 0 $X=563510 $Y=201805
X173 4 3 DCAPBWP7T $T=573320 241240 1 0 $X=573030 $Y=237030
X174 4 3 DCAPBWP7T $T=589000 209880 0 0 $X=588710 $Y=209645
X175 4 3 DCAPBWP7T $T=589560 170680 0 0 $X=589270 $Y=170445
X176 4 3 DCAPBWP7T $T=599080 225560 0 0 $X=598790 $Y=225325
X177 4 3 DCAPBWP7T $T=600200 162840 1 0 $X=599910 $Y=158630
X178 4 3 DCAPBWP7T $T=606920 170680 0 0 $X=606630 $Y=170445
X179 4 3 DCAPBWP7T $T=615320 217720 0 0 $X=615030 $Y=217485
X180 4 3 DCAPBWP7T $T=615320 233400 1 0 $X=615030 $Y=229190
X181 4 3 DCAPBWP7T $T=618120 202040 1 0 $X=617830 $Y=197830
X182 4 3 DCAPBWP7T $T=624840 241240 1 0 $X=624550 $Y=237030
X183 4 3 DCAPBWP7T $T=630440 178520 1 0 $X=630150 $Y=174310
X184 4 3 DCAPBWP7T $T=636600 241240 1 0 $X=636310 $Y=237030
X185 4 3 DCAPBWP7T $T=640520 225560 0 0 $X=640230 $Y=225325
X186 4 3 DCAPBWP7T $T=642200 170680 0 0 $X=641910 $Y=170445
X187 4 3 DCAPBWP7T $T=657320 178520 0 0 $X=657030 $Y=178285
X188 4 3 DCAPBWP7T $T=657320 209880 0 0 $X=657030 $Y=209645
X189 4 3 DCAPBWP7T $T=657320 225560 0 0 $X=657030 $Y=225325
X190 4 3 DCAPBWP7T $T=660120 170680 0 0 $X=659830 $Y=170445
X191 4 3 DCAPBWP7T $T=674680 202040 1 0 $X=674390 $Y=197830
X192 4 3 DCAPBWP7T $T=687000 225560 1 0 $X=686710 $Y=221350
X193 4 3 DCAPBWP7T $T=687560 241240 1 0 $X=687270 $Y=237030
X194 4 3 DCAPBWP7T $T=688680 194200 0 0 $X=688390 $Y=193965
X195 4 3 DCAPBWP7T $T=691480 186360 1 0 $X=691190 $Y=182150
X196 4 3 DCAPBWP7T $T=699320 178520 1 0 $X=699030 $Y=174310
X197 4 3 DCAPBWP7T $T=699320 202040 0 0 $X=699030 $Y=201805
X198 4 3 DCAPBWP7T $T=699320 209880 0 0 $X=699030 $Y=209645
X199 4 3 DCAPBWP7T $T=699320 241240 1 0 $X=699030 $Y=237030
X200 4 3 DCAPBWP7T $T=722280 194200 1 0 $X=721990 $Y=189990
X201 4 3 DCAPBWP7T $T=730680 225560 0 0 $X=730390 $Y=225325
X202 3 4 DCAP8BWP7T $T=450120 202040 0 0 $X=449830 $Y=201805
X203 3 4 DCAP8BWP7T $T=459080 202040 1 0 $X=458790 $Y=197830
X204 3 4 DCAP8BWP7T $T=463000 186360 0 0 $X=462710 $Y=186125
X205 3 4 DCAP8BWP7T $T=485960 162840 0 0 $X=485670 $Y=162605
X206 3 4 DCAP8BWP7T $T=485960 217720 1 0 $X=485670 $Y=213510
X207 3 4 DCAP8BWP7T $T=492120 170680 1 0 $X=491830 $Y=166470
X208 3 4 DCAP8BWP7T $T=492120 202040 1 0 $X=491830 $Y=197830
X209 3 4 DCAP8BWP7T $T=516760 178520 1 0 $X=516470 $Y=174310
X210 3 4 DCAP8BWP7T $T=526840 178520 1 0 $X=526550 $Y=174310
X211 3 4 DCAP8BWP7T $T=526840 241240 1 0 $X=526550 $Y=237030
X212 3 4 DCAP8BWP7T $T=527400 170680 0 0 $X=527110 $Y=170445
X213 3 4 DCAP8BWP7T $T=527400 225560 1 0 $X=527110 $Y=221350
X214 3 4 DCAP8BWP7T $T=527960 186360 0 0 $X=527670 $Y=186125
X215 3 4 DCAP8BWP7T $T=528520 209880 1 0 $X=528230 $Y=205670
X216 3 4 DCAP8BWP7T $T=528520 225560 0 0 $X=528230 $Y=225325
X217 3 4 DCAP8BWP7T $T=534120 202040 1 0 $X=533830 $Y=197830
X218 3 4 DCAP8BWP7T $T=552040 194200 1 0 $X=551750 $Y=189990
X219 3 4 DCAP8BWP7T $T=552040 217720 0 0 $X=551750 $Y=217485
X220 3 4 DCAP8BWP7T $T=569400 202040 1 0 $X=569110 $Y=197830
X221 3 4 DCAP8BWP7T $T=570520 186360 1 0 $X=570230 $Y=182150
X222 3 4 DCAP8BWP7T $T=576120 233400 0 0 $X=575830 $Y=233165
X223 3 4 DCAP8BWP7T $T=585080 170680 0 0 $X=584790 $Y=170445
X224 3 4 DCAP8BWP7T $T=585080 202040 1 0 $X=584790 $Y=197830
X225 3 4 DCAP8BWP7T $T=585080 209880 1 0 $X=584790 $Y=205670
X226 3 4 DCAP8BWP7T $T=594040 241240 1 0 $X=593750 $Y=237030
X227 3 4 DCAP8BWP7T $T=597960 194200 1 0 $X=597670 $Y=189990
X228 3 4 DCAP8BWP7T $T=602440 170680 0 0 $X=602150 $Y=170445
X229 3 4 DCAP8BWP7T $T=611400 233400 0 0 $X=611110 $Y=233165
X230 3 4 DCAP8BWP7T $T=611960 186360 1 0 $X=611670 $Y=182150
X231 3 4 DCAP8BWP7T $T=611960 209880 1 0 $X=611670 $Y=205670
X232 3 4 DCAP8BWP7T $T=612520 194200 1 0 $X=612230 $Y=189990
X233 3 4 DCAP8BWP7T $T=625960 178520 1 0 $X=625670 $Y=174310
X234 3 4 DCAP8BWP7T $T=627080 186360 0 0 $X=626790 $Y=186125
X235 3 4 DCAP8BWP7T $T=645000 202040 0 0 $X=644710 $Y=201805
X236 3 4 DCAP8BWP7T $T=652840 225560 0 0 $X=652550 $Y=225325
X237 3 4 DCAP8BWP7T $T=653960 162840 1 0 $X=653670 $Y=158630
X238 3 4 DCAP8BWP7T $T=654520 186360 0 0 $X=654230 $Y=186125
X239 3 4 DCAP8BWP7T $T=654520 233400 0 0 $X=654230 $Y=233165
X240 3 4 DCAP8BWP7T $T=660120 241240 1 0 $X=659830 $Y=237030
X241 3 4 DCAP8BWP7T $T=672440 202040 0 0 $X=672150 $Y=201805
X242 3 4 DCAP8BWP7T $T=687000 186360 1 0 $X=686710 $Y=182150
X243 3 4 DCAP8BWP7T $T=695960 170680 0 0 $X=695670 $Y=170445
X244 3 4 DCAP8BWP7T $T=695960 194200 1 0 $X=695670 $Y=189990
X245 3 4 DCAP8BWP7T $T=695960 202040 1 0 $X=695670 $Y=197830
X246 3 4 DCAP8BWP7T $T=696520 217720 0 0 $X=696230 $Y=217485
X247 3 4 DCAP8BWP7T $T=696520 233400 1 0 $X=696230 $Y=229190
X248 3 4 DCAP8BWP7T $T=702120 170680 1 0 $X=701830 $Y=166470
X249 3 4 DCAP8BWP7T $T=702120 209880 1 0 $X=701830 $Y=205670
X250 3 4 DCAP8BWP7T $T=717800 194200 1 0 $X=717510 $Y=189990
X251 3 4 DCAP8BWP7T $T=729560 170680 1 0 $X=729270 $Y=166470
X252 3 4 DCAP8BWP7T $T=737400 209880 1 0 $X=737110 $Y=205670
X253 3 4 DCAP8BWP7T $T=738520 170680 1 0 $X=738230 $Y=166470
X254 3 4 DCAP8BWP7T $T=738520 186360 1 0 $X=738230 $Y=182150
X255 3 4 DCAP8BWP7T $T=738520 194200 0 0 $X=738230 $Y=193965
X256 3 4 DCAP8BWP7T $T=738520 217720 1 0 $X=738230 $Y=213510
X257 3 4 DCAP8BWP7T $T=738520 225560 1 0 $X=738230 $Y=221350
X258 3 4 DCAP8BWP7T $T=738520 241240 1 0 $X=738230 $Y=237030
X259 3 4 DCAP4BWP7T $T=473080 209880 0 0 $X=472790 $Y=209645
X260 3 4 DCAP4BWP7T $T=473640 162840 1 0 $X=473350 $Y=158630
X261 3 4 DCAP4BWP7T $T=495480 170680 0 0 $X=495190 $Y=170445
X262 3 4 DCAP4BWP7T $T=501080 217720 1 0 $X=500790 $Y=213510
X263 3 4 DCAP4BWP7T $T=541400 225560 1 0 $X=541110 $Y=221350
X264 3 4 DCAP4BWP7T $T=572200 233400 0 0 $X=571910 $Y=233165
X265 3 4 DCAP4BWP7T $T=572760 155000 0 0 $X=572470 $Y=154765
X266 3 4 DCAP4BWP7T $T=585080 186360 1 0 $X=584790 $Y=182150
X267 3 4 DCAP4BWP7T $T=614200 186360 0 0 $X=613910 $Y=186125
X268 3 4 DCAP4BWP7T $T=614760 194200 0 0 $X=614470 $Y=193965
X269 3 4 DCAP4BWP7T $T=614760 202040 0 0 $X=614470 $Y=201805
X270 3 4 DCAP4BWP7T $T=614760 217720 1 0 $X=614470 $Y=213510
X271 3 4 DCAP4BWP7T $T=625400 186360 1 0 $X=625110 $Y=182150
X272 3 4 DCAP4BWP7T $T=656200 209880 1 0 $X=655910 $Y=205670
X273 3 4 DCAP4BWP7T $T=656200 225560 1 0 $X=655910 $Y=221350
X274 3 4 DCAP4BWP7T $T=656200 233400 1 0 $X=655910 $Y=229190
X275 3 4 DCAP4BWP7T $T=656760 194200 0 0 $X=656470 $Y=193965
X276 3 4 DCAP4BWP7T $T=656760 202040 1 0 $X=656470 $Y=197830
X277 3 4 DCAP4BWP7T $T=664040 225560 0 0 $X=663750 $Y=225325
X278 3 4 DCAP4BWP7T $T=669640 170680 0 0 $X=669350 $Y=170445
X279 3 4 DCAP4BWP7T $T=685880 217720 0 0 $X=685590 $Y=217485
X280 3 4 DCAP4BWP7T $T=691480 217720 0 0 $X=691190 $Y=217485
X281 3 4 DCAP4BWP7T $T=698200 178520 0 0 $X=697910 $Y=178285
X282 3 4 DCAP4BWP7T $T=698200 217720 1 0 $X=697910 $Y=213510
X283 3 4 DCAP4BWP7T $T=702120 233400 0 0 $X=701830 $Y=233165
X284 3 4 DCAP4BWP7T $T=717800 225560 0 0 $X=717510 $Y=225325
X285 3 4 DCAP4BWP7T $T=725640 186360 0 0 $X=725350 $Y=186125
X286 3 4 DCAP4BWP7T $T=740200 202040 1 0 $X=739910 $Y=197830
X287 3 4 DCAP4BWP7T $T=740200 209880 0 0 $X=739910 $Y=209645
X288 3 4 DCAP4BWP7T $T=740200 217720 0 0 $X=739910 $Y=217485
X289 3 4 ICV_40 $T=450120 155000 0 0 $X=449830 $Y=154765
X290 3 4 ICV_40 $T=474760 225560 0 0 $X=474470 $Y=225325
X291 3 4 ICV_40 $T=483160 202040 0 0 $X=482870 $Y=201805
X292 3 4 ICV_40 $T=483720 194200 1 0 $X=483430 $Y=189990
X293 3 4 ICV_40 $T=484280 233400 1 0 $X=483990 $Y=229190
X294 3 4 ICV_40 $T=492120 178520 0 0 $X=491830 $Y=178285
X295 3 4 ICV_40 $T=492120 225560 0 0 $X=491830 $Y=225325
X296 3 4 ICV_40 $T=501080 202040 1 0 $X=500790 $Y=197830
X297 3 4 ICV_40 $T=501080 225560 1 0 $X=500790 $Y=221350
X298 3 4 ICV_40 $T=510040 209880 0 0 $X=509750 $Y=209645
X299 3 4 ICV_40 $T=524600 170680 1 0 $X=524310 $Y=166470
X300 3 4 ICV_40 $T=524600 194200 1 0 $X=524310 $Y=189990
X301 3 4 ICV_40 $T=524600 233400 1 0 $X=524310 $Y=229190
X302 3 4 ICV_40 $T=534120 241240 1 0 $X=533830 $Y=237030
X303 3 4 ICV_40 $T=552040 155000 0 0 $X=551750 $Y=154765
X304 3 4 ICV_40 $T=552040 178520 0 0 $X=551750 $Y=178285
X305 3 4 ICV_40 $T=552040 233400 1 0 $X=551750 $Y=229190
X306 3 4 ICV_40 $T=557080 202040 0 0 $X=556790 $Y=201805
X307 3 4 ICV_40 $T=566600 241240 1 0 $X=566310 $Y=237030
X308 3 4 ICV_40 $T=567160 178520 1 0 $X=566870 $Y=174310
X309 3 4 ICV_40 $T=567720 170680 1 0 $X=567430 $Y=166470
X310 3 4 ICV_40 $T=568280 194200 1 0 $X=567990 $Y=189990
X311 3 4 ICV_40 $T=568280 202040 0 0 $X=567990 $Y=201805
X312 3 4 ICV_40 $T=582280 209880 0 0 $X=581990 $Y=209645
X313 3 4 ICV_40 $T=592360 225560 0 0 $X=592070 $Y=225325
X314 3 4 ICV_40 $T=596280 202040 0 0 $X=595990 $Y=201805
X315 3 4 ICV_40 $T=609720 162840 0 0 $X=609430 $Y=162605
X316 3 4 ICV_40 $T=618120 194200 0 0 $X=617830 $Y=193965
X317 3 4 ICV_40 $T=618120 241240 1 0 $X=617830 $Y=237030
X318 3 4 ICV_40 $T=627080 233400 1 0 $X=626790 $Y=229190
X319 3 4 ICV_40 $T=635480 170680 0 0 $X=635190 $Y=170445
X320 3 4 ICV_40 $T=638280 233400 0 0 $X=637990 $Y=233165
X321 3 4 ICV_40 $T=651720 178520 1 0 $X=651430 $Y=174310
X322 3 4 ICV_40 $T=652280 170680 1 0 $X=651990 $Y=166470
X323 3 4 ICV_40 $T=652280 202040 0 0 $X=651990 $Y=201805
X324 3 4 ICV_40 $T=660120 170680 1 0 $X=659830 $Y=166470
X325 3 4 ICV_40 $T=660120 186360 0 0 $X=659830 $Y=186125
X326 3 4 ICV_40 $T=692600 178520 1 0 $X=692310 $Y=174310
X327 3 4 ICV_40 $T=692600 209880 0 0 $X=692310 $Y=209645
X328 3 4 ICV_40 $T=692600 241240 1 0 $X=692310 $Y=237030
X329 3 4 ICV_40 $T=702120 225560 0 0 $X=701830 $Y=225325
X330 3 4 ICV_40 $T=720040 202040 0 0 $X=719750 $Y=201805
X331 3 4 ICV_40 $T=720600 178520 1 0 $X=720310 $Y=174310
X332 3 4 ICV_40 $T=728440 225560 1 0 $X=728150 $Y=221350
X333 3 4 ICV_40 $T=735160 162840 0 0 $X=734870 $Y=162605
X334 3 4 ICV_40 $T=735160 225560 0 0 $X=734870 $Y=225325
X335 3 4 ICV_40 $T=736280 194200 1 0 $X=735990 $Y=189990
X336 3 4 ICV_40 $T=736280 233400 0 0 $X=735990 $Y=233165
X337 4 3 DCAP64BWP7T $T=621480 178520 0 0 $X=621190 $Y=178285
X377 3 4 ICV_47 $T=450120 170680 1 0 $X=449830 $Y=166470
X378 3 4 ICV_47 $T=450120 178520 0 0 $X=449830 $Y=178285
X379 3 4 ICV_47 $T=450120 194200 0 0 $X=449830 $Y=193965
X380 3 4 ICV_47 $T=450120 225560 1 0 $X=449830 $Y=221350
X381 3 4 ICV_47 $T=450120 233400 0 0 $X=449830 $Y=233165
X382 3 4 ICV_47 $T=492120 155000 0 0 $X=491830 $Y=154765
X383 3 4 ICV_47 $T=492120 162840 0 0 $X=491830 $Y=162605
X384 3 4 ICV_47 $T=492120 202040 0 0 $X=491830 $Y=201805
X385 3 4 ICV_47 $T=576120 155000 0 0 $X=575830 $Y=154765
X386 3 4 ICV_47 $T=576120 178520 0 0 $X=575830 $Y=178285
X387 3 4 ICV_47 $T=618120 155000 0 0 $X=617830 $Y=154765
X388 3 4 ICV_47 $T=618120 162840 0 0 $X=617830 $Y=162605
X389 3 4 ICV_47 $T=660120 155000 0 0 $X=659830 $Y=154765
X390 3 4 ICV_47 $T=660120 162840 0 0 $X=659830 $Y=162605
X391 3 4 ICV_47 $T=702120 155000 0 0 $X=701830 $Y=154765
X392 3 4 ICV_47 $T=702120 178520 0 0 $X=701830 $Y=178285
X393 3 4 ICV_47 $T=702120 233400 1 0 $X=701830 $Y=229190
X394 4 3 DCAP32BWP7T $T=450120 162840 0 0 $X=449830 $Y=162605
X395 4 3 DCAP32BWP7T $T=450120 209880 1 0 $X=449830 $Y=205670
X396 4 3 DCAP32BWP7T $T=465240 202040 0 0 $X=464950 $Y=201805
X397 4 3 DCAP32BWP7T $T=465800 194200 1 0 $X=465510 $Y=189990
X398 4 3 DCAP32BWP7T $T=472520 155000 0 0 $X=472230 $Y=154765
X399 4 3 DCAP32BWP7T $T=492120 209880 0 0 $X=491830 $Y=209645
X400 4 3 DCAP32BWP7T $T=504440 194200 0 0 $X=504150 $Y=193965
X401 4 3 DCAP32BWP7T $T=505560 217720 0 0 $X=505270 $Y=217485
X402 4 3 DCAP32BWP7T $T=534120 155000 0 0 $X=533830 $Y=154765
X403 4 3 DCAP32BWP7T $T=534120 178520 0 0 $X=533830 $Y=178285
X404 4 3 DCAP32BWP7T $T=534120 194200 1 0 $X=533830 $Y=189990
X405 4 3 DCAP32BWP7T $T=534120 217720 0 0 $X=533830 $Y=217485
X406 4 3 DCAP32BWP7T $T=542520 202040 1 0 $X=542230 $Y=197830
X407 4 3 DCAP32BWP7T $T=545320 194200 0 0 $X=545030 $Y=193965
X408 4 3 DCAP32BWP7T $T=554280 233400 0 0 $X=553990 $Y=233165
X409 4 3 DCAP32BWP7T $T=556520 186360 0 0 $X=556230 $Y=186125
X410 4 3 DCAP32BWP7T $T=557080 217720 1 0 $X=556790 $Y=213510
X411 4 3 DCAP32BWP7T $T=557080 225560 0 0 $X=556790 $Y=225325
X412 4 3 DCAP32BWP7T $T=576120 162840 0 0 $X=575830 $Y=162605
X413 4 3 DCAP32BWP7T $T=576120 194200 1 0 $X=575830 $Y=189990
X414 4 3 DCAP32BWP7T $T=584520 233400 0 0 $X=584230 $Y=233165
X415 4 3 DCAP32BWP7T $T=587880 217720 1 0 $X=587590 $Y=213510
X416 4 3 DCAP32BWP7T $T=597400 217720 0 0 $X=597110 $Y=217485
X417 4 3 DCAP32BWP7T $T=618120 202040 0 0 $X=617830 $Y=201805
X418 4 3 DCAP32BWP7T $T=618120 217720 0 0 $X=617830 $Y=217485
X419 4 3 DCAP32BWP7T $T=625400 170680 1 0 $X=625110 $Y=166470
X420 4 3 DCAP32BWP7T $T=626520 194200 1 0 $X=626230 $Y=189990
X421 4 3 DCAP32BWP7T $T=629320 225560 1 0 $X=629030 $Y=221350
X422 4 3 DCAP32BWP7T $T=637720 217720 1 0 $X=637430 $Y=213510
X423 4 3 DCAP32BWP7T $T=641080 241240 1 0 $X=640790 $Y=237030
X424 4 3 DCAP32BWP7T $T=660120 178520 1 0 $X=659830 $Y=174310
X425 4 3 DCAP32BWP7T $T=660120 186360 1 0 $X=659830 $Y=182150
X426 4 3 DCAP32BWP7T $T=660120 225560 1 0 $X=659830 $Y=221350
X427 4 3 DCAP32BWP7T $T=660120 233400 1 0 $X=659830 $Y=229190
X428 4 3 DCAP32BWP7T $T=664040 209880 0 0 $X=663750 $Y=209645
X429 4 3 DCAP32BWP7T $T=671320 178520 0 0 $X=671030 $Y=178285
X430 4 3 DCAP32BWP7T $T=680280 217720 1 0 $X=679990 $Y=213510
X431 4 3 DCAP32BWP7T $T=682520 233400 0 0 $X=682230 $Y=233165
X432 4 3 DCAP32BWP7T $T=702120 162840 0 0 $X=701830 $Y=162605
X433 4 3 DCAP32BWP7T $T=702120 194200 0 0 $X=701830 $Y=193965
X434 4 3 DCAP32BWP7T $T=702120 202040 0 0 $X=701830 $Y=201805
X435 4 3 DCAP32BWP7T $T=702120 217720 1 0 $X=701830 $Y=213510
X436 4 3 DCAP32BWP7T $T=710520 209880 1 0 $X=710230 $Y=205670
X437 4 3 DCAP32BWP7T $T=722280 202040 1 0 $X=721990 $Y=197830
X554 52 3 37 57 4 ND2D1BWP7T $T=564360 241240 1 0 $X=564070 $Y=237030
X555 98 3 306 99 4 ND2D1BWP7T $T=692040 233400 1 0 $X=691750 $Y=229190
X556 98 3 101 57 4 ND2D1BWP7T $T=694280 233400 1 0 $X=693990 $Y=229190
X557 7 8 11 114 3 4 OAI21D0BWP7T $T=450680 241240 1 0 $X=450390 $Y=237030
X558 6 115 14 113 3 4 OAI21D0BWP7T $T=452920 186360 1 0 $X=452630 $Y=182150
X559 118 120 21 128 3 4 OAI21D0BWP7T $T=458520 155000 0 0 $X=458230 $Y=154765
X560 118 121 23 146 3 4 OAI21D0BWP7T $T=459640 186360 1 0 $X=459350 $Y=182150
X561 118 124 24 123 3 4 OAI21D0BWP7T $T=461880 170680 0 0 $X=461590 $Y=170445
X562 118 117 28 127 3 4 OAI21D0BWP7T $T=469720 217720 1 180 $X=466630 $Y=217485
X563 118 129 14 132 3 4 OAI21D0BWP7T $T=468600 209880 1 0 $X=468310 $Y=205670
X564 30 133 11 140 3 4 OAI21D0BWP7T $T=472520 233400 1 0 $X=472230 $Y=229190
X565 118 126 33 137 3 4 OAI21D0BWP7T $T=474760 217720 0 0 $X=474470 $Y=217485
X566 30 131 34 139 3 4 OAI21D0BWP7T $T=478120 241240 1 0 $X=477830 $Y=237030
X567 118 143 37 135 3 4 OAI21D0BWP7T $T=485960 162840 1 180 $X=482870 $Y=162605
X568 41 144 21 150 3 4 OAI21D0BWP7T $T=492680 170680 0 0 $X=492390 $Y=170445
X569 41 152 24 157 3 4 OAI21D0BWP7T $T=497720 170680 0 0 $X=497430 $Y=170445
X570 118 145 43 142 3 4 OAI21D0BWP7T $T=498280 202040 1 0 $X=497990 $Y=197830
X571 28 158 44 178 3 4 OAI21D0BWP7T $T=498840 225560 0 0 $X=498550 $Y=225325
X572 41 153 23 162 3 4 OAI21D0BWP7T $T=499960 178520 0 0 $X=499670 $Y=178285
X573 41 151 28 156 3 4 OAI21D0BWP7T $T=503320 217720 1 0 $X=503030 $Y=213510
X574 41 154 14 163 3 4 OAI21D0BWP7T $T=507800 209880 1 0 $X=507510 $Y=205670
X575 41 155 33 164 3 4 OAI21D0BWP7T $T=509480 225560 1 0 $X=509190 $Y=221350
X576 41 159 37 166 3 4 OAI21D0BWP7T $T=510600 178520 1 0 $X=510310 $Y=174310
X577 11 48 47 46 3 4 OAI21D0BWP7T $T=517880 241240 0 180 $X=514790 $Y=237030
X578 21 179 44 169 3 4 OAI21D0BWP7T $T=524600 170680 0 180 $X=521510 $Y=166470
X579 41 167 43 171 3 4 OAI21D0BWP7T $T=524600 194200 0 180 $X=521510 $Y=189990
X580 33 182 44 184 3 4 OAI21D0BWP7T $T=524600 225560 1 0 $X=524310 $Y=221350
X581 37 186 44 190 3 4 OAI21D0BWP7T $T=534680 170680 1 0 $X=534390 $Y=166470
X582 14 183 44 191 3 4 OAI21D0BWP7T $T=534680 209880 1 0 $X=534390 $Y=205670
X583 23 185 44 187 3 4 OAI21D0BWP7T $T=535240 186360 1 0 $X=534950 $Y=182150
X584 44 194 43 188 3 4 OAI21D0BWP7T $T=542520 202040 0 180 $X=539430 $Y=197830
X585 53 209 56 212 3 4 OAI21D0BWP7T $T=564360 178520 1 0 $X=564070 $Y=174310
X586 54 210 53 211 3 4 OAI21D0BWP7T $T=564360 194200 0 0 $X=564070 $Y=193965
X587 55 207 53 213 3 4 OAI21D0BWP7T $T=565480 202040 0 0 $X=565190 $Y=201805
X588 24 204 44 196 3 4 OAI21D0BWP7T $T=570520 162840 0 180 $X=567430 $Y=158630
X589 54 205 60 217 3 4 OAI21D0BWP7T $T=576680 217720 0 0 $X=576390 $Y=217485
X590 55 208 60 218 3 4 OAI21D0BWP7T $T=576680 233400 1 0 $X=576390 $Y=229190
X591 61 63 56 64 3 4 OAI21D0BWP7T $T=581720 233400 0 0 $X=581430 $Y=233165
X592 60 216 56 223 3 4 OAI21D0BWP7T $T=585080 217720 1 0 $X=584790 $Y=213510
X593 55 224 65 236 3 4 OAI21D0BWP7T $T=588440 225560 1 0 $X=588150 $Y=221350
X594 54 230 65 227 3 4 OAI21D0BWP7T $T=593480 202040 0 180 $X=590390 $Y=197830
X595 65 225 56 234 3 4 OAI21D0BWP7T $T=595160 194200 1 0 $X=594870 $Y=189990
X596 54 239 68 241 3 4 OAI21D0BWP7T $T=603000 202040 0 0 $X=602710 $Y=201805
X597 68 240 56 244 3 4 OAI21D0BWP7T $T=603560 194200 1 0 $X=603270 $Y=189990
X598 55 242 68 243 3 4 OAI21D0BWP7T $T=605240 225560 1 0 $X=604950 $Y=221350
X599 71 247 56 250 3 4 OAI21D0BWP7T $T=618680 178520 0 0 $X=618390 $Y=178285
X600 54 248 71 253 3 4 OAI21D0BWP7T $T=619800 202040 1 0 $X=619510 $Y=197830
X601 55 254 71 265 3 4 OAI21D0BWP7T $T=623160 217720 1 0 $X=622870 $Y=213510
X602 73 261 56 252 3 4 OAI21D0BWP7T $T=630440 186360 0 180 $X=627350 $Y=182150
X603 54 266 73 257 3 4 OAI21D0BWP7T $T=633800 186360 0 0 $X=633510 $Y=186125
X604 55 267 73 260 3 4 OAI21D0BWP7T $T=635480 233400 1 0 $X=635190 $Y=229190
X605 82 272 83 274 3 4 OAI21D0BWP7T $T=645000 233400 0 0 $X=644710 $Y=233165
X606 84 273 85 276 3 4 OAI21D0BWP7T $T=647240 186360 1 0 $X=646950 $Y=182150
X607 86 269 84 281 3 4 OAI21D0BWP7T $T=649480 202040 0 0 $X=649190 $Y=201805
X608 89 286 84 283 3 4 OAI21D0BWP7T $T=664040 194200 1 180 $X=660950 $Y=193965
X609 90 270 84 288 3 4 OAI21D0BWP7T $T=661240 209880 0 0 $X=660950 $Y=209645
X610 84 285 88 278 3 4 OAI21D0BWP7T $T=661240 225560 0 0 $X=660950 $Y=225325
X611 85 302 83 293 3 4 OAI21D0BWP7T $T=666840 170680 1 0 $X=666550 $Y=166470
X612 86 294 83 291 3 4 OAI21D0BWP7T $T=670200 186360 1 180 $X=667110 $Y=186125
X613 83 303 88 287 3 4 OAI21D0BWP7T $T=676920 217720 1 180 $X=673830 $Y=217485
X614 89 304 83 301 3 4 OAI21D0BWP7T $T=678040 170680 1 180 $X=674950 $Y=170445
X615 90 305 83 296 3 4 OAI21D0BWP7T $T=679720 202040 1 180 $X=676630 $Y=201805
X616 82 299 306 292 3 4 OAI21D0BWP7T $T=682520 233400 1 180 $X=679430 $Y=233165
X617 89 310 306 312 3 4 OAI21D0BWP7T $T=684200 170680 0 0 $X=683910 $Y=170445
X618 306 311 88 313 3 4 OAI21D0BWP7T $T=691480 225560 0 180 $X=688390 $Y=221350
X619 90 314 306 316 3 4 OAI21D0BWP7T $T=689240 209880 1 0 $X=688950 $Y=205670
X620 86 309 306 319 3 4 OAI21D0BWP7T $T=690360 194200 0 0 $X=690070 $Y=193965
X621 306 318 85 321 3 4 OAI21D0BWP7T $T=692600 170680 1 0 $X=692310 $Y=166470
X622 90 320 100 322 3 4 OAI21D0BWP7T $T=693720 217720 0 0 $X=693430 $Y=217485
X623 86 324 100 325 3 4 OAI21D0BWP7T $T=707720 209880 1 0 $X=707430 $Y=205670
X624 89 336 100 335 3 4 OAI21D0BWP7T $T=716680 186360 1 180 $X=713590 $Y=186125
X625 100 338 85 351 3 4 OAI21D0BWP7T $T=721720 170680 0 0 $X=721430 $Y=170445
X626 90 340 101 332 3 4 OAI21D0BWP7T $T=724520 233400 0 0 $X=724230 $Y=233165
X627 86 345 101 328 3 4 OAI21D0BWP7T $T=732360 225560 0 0 $X=732070 $Y=225325
X628 106 107 85 348 3 4 OAI21D0BWP7T $T=732360 241240 1 0 $X=732070 $Y=237030
X629 101 350 85 341 3 4 OAI21D0BWP7T $T=738520 217720 0 180 $X=735430 $Y=213510
X630 89 346 101 347 3 4 OAI21D0BWP7T $T=738520 225560 0 180 $X=735430 $Y=221350
X662 3 4 DCAP16BWP7T $T=454040 186360 0 0 $X=453750 $Y=186125
X663 3 4 DCAP16BWP7T $T=462440 233400 1 0 $X=462150 $Y=229190
X664 3 4 DCAP16BWP7T $T=464680 162840 1 0 $X=464390 $Y=158630
X665 3 4 DCAP16BWP7T $T=469720 217720 1 0 $X=469430 $Y=213510
X666 3 4 DCAP16BWP7T $T=478120 170680 0 0 $X=477830 $Y=170445
X667 3 4 DCAP16BWP7T $T=481480 217720 0 0 $X=481190 $Y=217485
X668 3 4 DCAP16BWP7T $T=492120 194200 1 0 $X=491830 $Y=189990
X669 3 4 DCAP16BWP7T $T=492120 217720 1 0 $X=491830 $Y=213510
X670 3 4 DCAP16BWP7T $T=492120 225560 1 0 $X=491830 $Y=221350
X671 3 4 DCAP16BWP7T $T=503320 233400 0 0 $X=503030 $Y=233165
X672 3 4 DCAP16BWP7T $T=515640 233400 1 0 $X=515350 $Y=229190
X673 3 4 DCAP16BWP7T $T=519560 209880 1 0 $X=519270 $Y=205670
X674 3 4 DCAP16BWP7T $T=520680 178520 0 0 $X=520390 $Y=178285
X675 3 4 DCAP16BWP7T $T=522360 194200 0 0 $X=522070 $Y=193965
X676 3 4 DCAP16BWP7T $T=523480 217720 0 0 $X=523190 $Y=217485
X677 3 4 DCAP16BWP7T $T=534120 162840 0 0 $X=533830 $Y=162605
X678 3 4 DCAP16BWP7T $T=534120 186360 0 0 $X=533830 $Y=186125
X679 3 4 DCAP16BWP7T $T=538600 233400 0 0 $X=538310 $Y=233165
X680 3 4 DCAP16BWP7T $T=543080 233400 1 0 $X=542790 $Y=229190
X681 3 4 DCAP16BWP7T $T=547000 241240 1 0 $X=546710 $Y=237030
X682 3 4 DCAP16BWP7T $T=553720 178520 1 0 $X=553430 $Y=174310
X683 3 4 DCAP16BWP7T $T=557640 162840 1 0 $X=557350 $Y=158630
X684 3 4 DCAP16BWP7T $T=560440 202040 1 0 $X=560150 $Y=197830
X685 3 4 DCAP16BWP7T $T=562680 170680 0 0 $X=562390 $Y=170445
X686 3 4 DCAP16BWP7T $T=563800 155000 0 0 $X=563510 $Y=154765
X687 3 4 DCAP16BWP7T $T=565480 225560 1 0 $X=565190 $Y=221350
X688 3 4 DCAP16BWP7T $T=566040 162840 0 0 $X=565750 $Y=162605
X689 3 4 DCAP16BWP7T $T=583400 225560 0 0 $X=583110 $Y=225325
X690 3 4 DCAP16BWP7T $T=600760 162840 0 0 $X=600470 $Y=162605
X691 3 4 DCAP16BWP7T $T=602440 233400 0 0 $X=602150 $Y=233165
X692 3 4 DCAP16BWP7T $T=605240 186360 0 0 $X=604950 $Y=186125
X693 3 4 DCAP16BWP7T $T=605800 202040 0 0 $X=605510 $Y=201805
X694 3 4 DCAP16BWP7T $T=605800 217720 1 0 $X=605510 $Y=213510
X695 3 4 DCAP16BWP7T $T=608040 225560 1 0 $X=607750 $Y=221350
X696 3 4 DCAP16BWP7T $T=618120 170680 0 0 $X=617830 $Y=170445
X697 3 4 DCAP16BWP7T $T=618120 186360 0 0 $X=617830 $Y=186125
X698 3 4 DCAP16BWP7T $T=629320 233400 0 0 $X=629030 $Y=233165
X699 3 4 DCAP16BWP7T $T=636040 202040 0 0 $X=635750 $Y=201805
X700 3 4 DCAP16BWP7T $T=636040 217720 0 0 $X=635750 $Y=217485
X701 3 4 DCAP16BWP7T $T=642760 178520 1 0 $X=642470 $Y=174310
X702 3 4 DCAP16BWP7T $T=643320 170680 1 0 $X=643030 $Y=166470
X703 3 4 DCAP16BWP7T $T=644440 194200 1 0 $X=644150 $Y=189990
X704 3 4 DCAP16BWP7T $T=647240 209880 1 0 $X=646950 $Y=205670
X705 3 4 DCAP16BWP7T $T=647240 225560 1 0 $X=646950 $Y=221350
X706 3 4 DCAP16BWP7T $T=647800 194200 0 0 $X=647510 $Y=193965
X707 3 4 DCAP16BWP7T $T=650040 186360 1 0 $X=649750 $Y=182150
X708 3 4 DCAP16BWP7T $T=676920 217720 0 0 $X=676630 $Y=217485
X709 3 4 DCAP16BWP7T $T=678040 186360 1 0 $X=677750 $Y=182150
X710 3 4 DCAP16BWP7T $T=678040 225560 1 0 $X=677750 $Y=221350
X711 3 4 DCAP16BWP7T $T=678040 233400 1 0 $X=677750 $Y=229190
X712 3 4 DCAP16BWP7T $T=679720 202040 0 0 $X=679430 $Y=201805
X713 3 4 DCAP16BWP7T $T=687000 202040 1 0 $X=686710 $Y=197830
X714 3 4 DCAP16BWP7T $T=688680 225560 0 0 $X=688390 $Y=225325
X715 3 4 DCAP16BWP7T $T=689240 178520 0 0 $X=688950 $Y=178285
X716 3 4 DCAP16BWP7T $T=691480 225560 1 0 $X=691190 $Y=221350
X717 3 4 DCAP16BWP7T $T=692040 209880 1 0 $X=691750 $Y=205670
X718 3 4 DCAP16BWP7T $T=702120 170680 0 0 $X=701830 $Y=170445
X719 3 4 DCAP16BWP7T $T=708840 194200 1 0 $X=708550 $Y=189990
X720 3 4 DCAP16BWP7T $T=711640 178520 1 0 $X=711350 $Y=174310
X721 3 4 DCAP16BWP7T $T=716680 186360 0 0 $X=716390 $Y=186125
X722 3 4 DCAP16BWP7T $T=726200 162840 0 0 $X=725910 $Y=162605
X723 3 4 DCAP16BWP7T $T=727320 194200 1 0 $X=727030 $Y=189990
X724 3 4 DCAP16BWP7T $T=727320 233400 0 0 $X=727030 $Y=233165
X725 3 4 DCAP16BWP7T $T=728440 209880 1 0 $X=728150 $Y=205670
X726 3 4 DCAP16BWP7T $T=729560 186360 1 0 $X=729270 $Y=182150
X727 3 4 DCAP16BWP7T $T=731240 209880 0 0 $X=730950 $Y=209645
X821 17 19 3 4 5 DFQD0BWP7T $T=461320 170680 1 180 $X=450390 $Y=170445
X822 17 20 3 4 9 DFQD0BWP7T $T=462440 233400 0 180 $X=451510 $Y=229190
X823 17 120 3 4 2 DFQD0BWP7T $T=464680 162840 0 180 $X=453750 $Y=158630
X824 17 117 3 4 125 DFQD0BWP7T $T=454600 202040 0 0 $X=454310 $Y=201805
X825 17 115 3 4 13 DFQD0BWP7T $T=465800 194200 0 180 $X=454870 $Y=189990
X826 17 126 3 4 119 DFQD0BWP7T $T=469720 217720 0 180 $X=458790 $Y=213510
X827 17 124 3 4 25 DFQD0BWP7T $T=473640 178520 0 180 $X=462710 $Y=174310
X828 17 131 3 4 26 DFQD0BWP7T $T=474760 225560 1 180 $X=463830 $Y=225325
X829 17 133 3 4 122 DFQD0BWP7T $T=475320 241240 0 180 $X=464390 $Y=237030
X830 17 129 3 4 116 DFQD0BWP7T $T=475880 202040 0 180 $X=464950 $Y=197830
X831 17 121 3 4 27 DFQD0BWP7T $T=478120 186360 1 180 $X=467190 $Y=186125
X832 45 42 3 4 39 DFQD0BWP7T $T=503320 233400 1 180 $X=492390 $Y=233165
X833 45 152 3 4 130 DFQD0BWP7T $T=503880 162840 0 180 $X=492950 $Y=158630
X834 17 151 3 4 147 DFQD0BWP7T $T=493240 209880 1 0 $X=492950 $Y=205670
X835 45 154 3 4 138 DFQD0BWP7T $T=504440 194200 1 180 $X=493510 $Y=193965
X836 45 153 3 4 149 DFQD0BWP7T $T=505560 186360 0 180 $X=494630 $Y=182150
X837 45 155 3 4 141 DFQD0BWP7T $T=505560 217720 1 180 $X=494630 $Y=217485
X838 45 158 3 4 168 DFQD0BWP7T $T=505000 233400 1 0 $X=504710 $Y=229190
X839 45 159 3 4 136 DFQD0BWP7T $T=505560 162840 1 0 $X=505270 $Y=158630
X840 45 167 3 4 148 DFQD0BWP7T $T=516760 194200 0 180 $X=505830 $Y=189990
X841 45 177 3 4 170 DFQD0BWP7T $T=517880 186360 1 0 $X=517590 $Y=182150
X842 45 186 3 4 172 DFQD0BWP7T $T=534680 162840 1 0 $X=534390 $Y=158630
X843 45 194 3 4 176 DFQD0BWP7T $T=545320 194200 1 180 $X=534390 $Y=193965
X844 45 185 3 4 165 DFQD0BWP7T $T=556520 186360 1 180 $X=545590 $Y=186125
X845 45 199 3 4 195 DFQD0BWP7T $T=557080 202040 1 180 $X=546150 $Y=201805
X846 45 201 3 4 189 DFQD0BWP7T $T=557080 217720 0 180 $X=546150 $Y=213510
X847 45 197 3 4 193 DFQD0BWP7T $T=557080 225560 1 180 $X=546150 $Y=225325
X848 45 204 3 4 161 DFQD0BWP7T $T=557640 162840 0 180 $X=546710 $Y=158630
X849 45 206 3 4 200 DFQD0BWP7T $T=567720 170680 0 180 $X=556790 $Y=166470
X850 45 203 3 4 202 DFQD0BWP7T $T=568280 194200 0 180 $X=557350 $Y=189990
X851 45 205 3 4 214 DFQD0BWP7T $T=558200 217720 0 0 $X=557910 $Y=217485
X852 45 207 3 4 58 DFQD0BWP7T $T=558760 209880 1 0 $X=558470 $Y=205670
X853 45 208 3 4 59 DFQD0BWP7T $T=559320 233400 1 0 $X=559030 $Y=229190
X854 45 215 3 4 221 DFQD0BWP7T $T=576680 162840 1 0 $X=576390 $Y=158630
X855 45 209 3 4 222 DFQD0BWP7T $T=576680 178520 1 0 $X=576390 $Y=174310
X856 45 210 3 4 219 DFQD0BWP7T $T=576680 186360 0 0 $X=576390 $Y=186125
X857 45 216 3 4 220 DFQD0BWP7T $T=576680 202040 0 0 $X=576390 $Y=201805
X858 45 224 3 4 69 DFQD0BWP7T $T=586760 233400 1 0 $X=586470 $Y=229190
X859 45 225 3 4 233 DFQD0BWP7T $T=587320 186360 1 0 $X=587030 $Y=182150
X860 45 232 3 4 226 DFQD0BWP7T $T=600200 162840 0 180 $X=589270 $Y=158630
X861 45 231 3 4 228 DFQD0BWP7T $T=601320 209880 1 180 $X=590390 $Y=209645
X862 45 240 3 4 245 DFQD0BWP7T $T=601320 186360 1 0 $X=601030 $Y=182150
X863 45 235 3 4 237 DFQD0BWP7T $T=601880 162840 1 0 $X=601590 $Y=158630
X864 45 239 3 4 246 DFQD0BWP7T $T=601880 209880 0 0 $X=601590 $Y=209645
X865 45 249 3 4 251 DFQD0BWP7T $T=618680 162840 1 0 $X=618390 $Y=158630
X866 45 248 3 4 262 DFQD0BWP7T $T=618680 209880 1 0 $X=618390 $Y=205670
X867 45 72 3 4 74 DFQD0BWP7T $T=618680 233400 0 0 $X=618390 $Y=233165
X868 81 266 3 4 259 DFQD0BWP7T $T=640520 202040 0 180 $X=629590 $Y=197830
X869 81 267 3 4 76 DFQD0BWP7T $T=640520 225560 1 180 $X=629590 $Y=225325
X870 81 254 3 4 78 DFQD0BWP7T $T=641080 209880 1 180 $X=630150 $Y=209645
X871 81 264 3 4 258 DFQD0BWP7T $T=642760 162840 0 180 $X=631830 $Y=158630
X872 81 247 3 4 256 DFQD0BWP7T $T=642760 178520 0 180 $X=631830 $Y=174310
X873 81 261 3 4 255 DFQD0BWP7T $T=648360 186360 1 180 $X=637430 $Y=186125
X874 81 269 3 4 279 DFQD0BWP7T $T=641640 202040 1 0 $X=641350 $Y=197830
X875 81 270 3 4 275 DFQD0BWP7T $T=642200 209880 0 0 $X=641910 $Y=209645
X876 81 271 3 4 282 DFQD0BWP7T $T=643320 162840 1 0 $X=643030 $Y=158630
X877 81 273 3 4 277 DFQD0BWP7T $T=643880 170680 0 0 $X=643590 $Y=170445
X878 81 286 3 4 280 DFQD0BWP7T $T=671320 178520 1 180 $X=660390 $Y=178285
X879 81 285 3 4 87 DFQD0BWP7T $T=676920 225560 1 180 $X=665990 $Y=225325
X880 81 303 3 4 284 DFQD0BWP7T $T=680280 217720 0 180 $X=669350 $Y=213510
X881 81 294 3 4 300 DFQD0BWP7T $T=670200 186360 0 0 $X=669910 $Y=186125
X882 81 302 3 4 295 DFQD0BWP7T $T=670760 162840 1 0 $X=670470 $Y=158630
X883 81 305 3 4 289 DFQD0BWP7T $T=687000 202040 0 180 $X=676070 $Y=197830
X884 81 311 3 4 290 DFQD0BWP7T $T=688680 225560 1 180 $X=677750 $Y=225325
X885 81 304 3 4 298 DFQD0BWP7T $T=692600 178520 0 180 $X=681670 $Y=174310
X886 81 309 3 4 315 DFQD0BWP7T $T=681960 186360 0 0 $X=681670 $Y=186125
X887 81 314 3 4 307 DFQD0BWP7T $T=692600 209880 1 180 $X=681670 $Y=209645
X888 81 318 3 4 326 DFQD0BWP7T $T=702680 162840 1 0 $X=702390 $Y=158630
X889 81 320 3 4 317 DFQD0BWP7T $T=702680 209880 0 0 $X=702390 $Y=209645
X890 81 324 3 4 327 DFQD0BWP7T $T=703240 202040 1 0 $X=702950 $Y=197830
X891 81 102 3 4 95 DFQD0BWP7T $T=715000 233400 1 180 $X=704070 $Y=233165
X892 81 310 3 4 323 DFQD0BWP7T $T=716120 186360 0 180 $X=705190 $Y=182150
X893 81 329 3 4 334 DFQD0BWP7T $T=726760 162840 0 180 $X=715830 $Y=158630
X894 81 336 3 4 330 DFQD0BWP7T $T=729560 186360 0 180 $X=718630 $Y=182150
X895 81 345 3 4 331 DFQD0BWP7T $T=730680 225560 1 180 $X=719750 $Y=225325
X896 81 346 3 4 333 DFQD0BWP7T $T=731240 209880 1 180 $X=720310 $Y=209645
X897 81 272 3 4 268 DFQD1BWP7T $T=652840 225560 1 180 $X=641910 $Y=225325
X898 81 299 3 4 92 DFQD1BWP7T $T=675240 241240 0 180 $X=664310 $Y=237030
X899 268 80 3 4 BUFFD1P5BWP7T $T=641080 241240 0 180 $X=637990 $Y=237030
X900 222 56 4 221 3 29 212 AOI22D1BWP7T $T=595160 170680 1 180 $X=590950 $Y=170445
X901 170 180 4 3 180 177 21 MAOI22D0BWP7T $T=526840 178520 0 180 $X=522630 $Y=174310
X902 173 180 4 3 180 181 28 MAOI22D0BWP7T $T=534680 233400 0 0 $X=534390 $Y=233165
X903 198 180 4 3 180 192 23 MAOI22D0BWP7T $T=541960 178520 0 180 $X=537750 $Y=174310
X904 193 180 4 3 180 197 14 MAOI22D0BWP7T $T=539160 233400 1 0 $X=538870 $Y=229190
X905 195 180 4 3 180 199 43 MAOI22D0BWP7T $T=540840 209880 0 0 $X=540550 $Y=209645
X906 189 180 4 3 180 201 33 MAOI22D0BWP7T $T=543640 225560 1 0 $X=543350 $Y=221350
X907 202 180 4 3 180 203 37 MAOI22D0BWP7T $T=548680 186360 1 0 $X=548390 $Y=182150
X908 200 180 4 3 180 206 24 MAOI22D0BWP7T $T=563800 155000 1 180 $X=559590 $Y=154765
X909 221 62 4 3 62 215 53 MAOI22D0BWP7T $T=585080 170680 0 180 $X=580870 $Y=166470
X910 66 62 4 3 62 229 61 MAOI22D0BWP7T $T=594040 241240 0 180 $X=589830 $Y=237030
X911 228 62 4 3 62 231 60 MAOI22D0BWP7T $T=597400 217720 1 180 $X=593190 $Y=217485
X912 237 62 4 3 62 235 68 MAOI22D0BWP7T $T=600760 162840 1 180 $X=596550 $Y=162605
X913 226 62 4 3 62 232 65 MAOI22D0BWP7T $T=598520 170680 0 0 $X=598230 $Y=170445
X914 251 62 4 3 62 249 73 MAOI22D0BWP7T $T=621480 170680 1 0 $X=621190 $Y=166470
X915 258 62 4 3 62 264 71 MAOI22D0BWP7T $T=635480 170680 1 180 $X=631270 $Y=170445
X916 282 91 4 3 91 271 84 MAOI22D0BWP7T $T=664600 162840 0 180 $X=660390 $Y=158630
X917 297 91 4 3 91 308 83 MAOI22D0BWP7T $T=685880 162840 0 180 $X=681670 $Y=158630
X918 334 91 4 3 91 329 306 MAOI22D0BWP7T $T=711640 170680 0 180 $X=707430 $Y=166470
X919 342 91 4 3 91 339 100 MAOI22D0BWP7T $T=726200 162840 1 180 $X=721990 $Y=162605
X920 344 91 4 3 91 349 101 MAOI22D0BWP7T $T=734600 194200 0 0 $X=734310 $Y=193965
X921 6 113 10 13 116 4 3 AOI22D0BWP7T $T=450680 186360 0 0 $X=450390 $Y=186125
X922 6 12 10 15 125 4 3 AOI22D0BWP7T $T=451800 209880 0 0 $X=451510 $Y=209645
X923 6 16 10 18 119 4 3 AOI22D0BWP7T $T=454600 217720 0 0 $X=454310 $Y=217485
X924 7 114 10 22 122 4 3 AOI22D0BWP7T $T=457400 241240 1 0 $X=457110 $Y=237030
X925 118 123 29 25 130 4 3 AOI22D0BWP7T $T=468040 162840 0 0 $X=467750 $Y=162605
X926 118 128 29 2 134 4 3 AOI22D0BWP7T $T=469160 155000 0 0 $X=468870 $Y=154765
X927 118 135 29 31 136 4 3 AOI22D0BWP7T $T=474760 170680 0 0 $X=474470 $Y=170445
X928 118 132 29 116 138 4 3 AOI22D0BWP7T $T=475320 209880 0 0 $X=475030 $Y=209645
X929 118 137 10 119 141 4 3 AOI22D0BWP7T $T=478120 217720 0 0 $X=477830 $Y=217485
X930 30 140 10 122 36 4 3 AOI22D0BWP7T $T=480920 233400 1 0 $X=480630 $Y=229190
X931 118 142 29 32 148 4 3 AOI22D0BWP7T $T=481480 209880 1 0 $X=481190 $Y=205670
X932 118 127 10 125 147 4 3 AOI22D0BWP7T $T=482600 217720 1 0 $X=482310 $Y=213510
X933 30 139 10 26 40 4 3 AOI22D0BWP7T $T=482600 241240 1 0 $X=482310 $Y=237030
X934 118 146 29 27 149 4 3 AOI22D0BWP7T $T=483160 186360 0 0 $X=482870 $Y=186125
X935 41 150 29 134 160 4 3 AOI22D0BWP7T $T=498840 170680 1 0 $X=498550 $Y=166470
X936 41 157 29 130 161 4 3 AOI22D0BWP7T $T=506120 170680 0 0 $X=505830 $Y=170445
X937 41 162 29 149 165 4 3 AOI22D0BWP7T $T=509480 186360 1 0 $X=509190 $Y=182150
X938 41 163 29 138 174 4 3 AOI22D0BWP7T $T=509480 202040 1 0 $X=509190 $Y=197830
X939 41 156 29 147 168 4 3 AOI22D0BWP7T $T=510600 217720 1 0 $X=510310 $Y=213510
X940 41 166 29 136 172 4 3 AOI22D0BWP7T $T=513400 178520 1 0 $X=513110 $Y=174310
X941 44 169 29 160 170 4 3 AOI22D0BWP7T $T=513960 170680 1 0 $X=513670 $Y=166470
X942 41 164 29 141 175 4 3 AOI22D0BWP7T $T=515080 225560 1 0 $X=514790 $Y=221350
X943 41 171 29 148 176 4 3 AOI22D0BWP7T $T=516200 209880 1 0 $X=515910 $Y=205670
X944 44 178 29 168 173 4 3 AOI22D0BWP7T $T=523480 225560 0 180 $X=519830 $Y=221350
X945 44 184 29 175 189 4 3 AOI22D0BWP7T $T=534680 225560 1 0 $X=534390 $Y=221350
X946 44 188 29 176 195 4 3 AOI22D0BWP7T $T=536920 209880 0 0 $X=536630 $Y=209645
X947 44 187 29 165 198 4 3 AOI22D0BWP7T $T=538040 186360 1 0 $X=537750 $Y=182150
X948 44 191 29 174 193 4 3 AOI22D0BWP7T $T=538040 225560 1 0 $X=537750 $Y=221350
X949 44 196 29 161 200 4 3 AOI22D0BWP7T $T=541400 170680 0 0 $X=541110 $Y=170445
X950 44 190 29 172 202 4 3 AOI22D0BWP7T $T=544760 162840 0 0 $X=544470 $Y=162605
X951 55 213 29 58 219 4 3 AOI22D0BWP7T $T=578920 209880 0 0 $X=578630 $Y=209645
X952 55 218 29 59 214 4 3 AOI22D0BWP7T $T=583400 225560 1 180 $X=579750 $Y=225325
X953 54 217 29 214 220 4 3 AOI22D0BWP7T $T=580600 217720 0 0 $X=580310 $Y=217485
X954 54 211 29 219 222 4 3 AOI22D0BWP7T $T=581160 194200 0 0 $X=580870 $Y=193965
X955 56 223 29 220 228 4 3 AOI22D0BWP7T $T=590680 209880 1 0 $X=590390 $Y=205670
X956 54 227 67 238 233 4 3 AOI22D0BWP7T $T=593480 194200 0 0 $X=593190 $Y=193965
X957 55 236 67 69 238 4 3 AOI22D0BWP7T $T=598520 241240 1 0 $X=598230 $Y=237030
X958 56 234 67 233 226 4 3 AOI22D0BWP7T $T=608040 178520 0 180 $X=604390 $Y=174310
X959 56 244 67 245 237 4 3 AOI22D0BWP7T $T=608600 170680 0 0 $X=608310 $Y=170445
X960 54 241 67 246 245 4 3 AOI22D0BWP7T $T=609160 194200 1 0 $X=608870 $Y=189990
X961 55 243 67 70 246 4 3 AOI22D0BWP7T $T=618680 225560 1 0 $X=618390 $Y=221350
X962 56 252 67 255 251 4 3 AOI22D0BWP7T $T=622040 186360 1 0 $X=621750 $Y=182150
X963 56 250 67 256 258 4 3 AOI22D0BWP7T $T=622600 178520 1 0 $X=622310 $Y=174310
X964 54 257 67 259 255 4 3 AOI22D0BWP7T $T=623160 194200 1 0 $X=622870 $Y=189990
X965 55 260 67 76 259 4 3 AOI22D0BWP7T $T=625960 225560 1 0 $X=625670 $Y=221350
X966 54 253 67 262 256 4 3 AOI22D0BWP7T $T=626520 194200 0 0 $X=626230 $Y=193965
X967 56 77 67 75 74 4 3 AOI22D0BWP7T $T=629880 241240 0 180 $X=626230 $Y=237030
X968 55 265 67 78 262 4 3 AOI22D0BWP7T $T=634360 217720 1 0 $X=634070 $Y=213510
X969 88 278 67 87 275 4 3 AOI22D0BWP7T $T=652280 217720 1 180 $X=648630 $Y=217485
X970 89 283 67 280 277 4 3 AOI22D0BWP7T $T=654520 186360 1 180 $X=650870 $Y=186125
X971 284 274 80 67 82 4 3 AOI22D0BWP7T $T=654520 233400 1 180 $X=650870 $Y=233165
X972 85 276 67 277 282 4 3 AOI22D0BWP7T $T=665160 170680 1 180 $X=661510 $Y=170445
X973 86 281 67 279 280 4 3 AOI22D0BWP7T $T=665720 202040 0 180 $X=662070 $Y=197830
X974 88 287 67 284 289 4 3 AOI22D0BWP7T $T=662360 217720 0 0 $X=662070 $Y=217485
X975 90 288 67 275 279 4 3 AOI22D0BWP7T $T=666280 209880 0 180 $X=662630 $Y=205670
X976 290 292 92 67 82 4 3 AOI22D0BWP7T $T=667400 233400 1 180 $X=663750 $Y=233165
X977 85 293 67 295 297 4 3 AOI22D0BWP7T $T=667400 162840 1 0 $X=667110 $Y=158630
X978 86 291 67 300 298 4 3 AOI22D0BWP7T $T=667400 194200 0 0 $X=667110 $Y=193965
X979 90 296 67 289 300 4 3 AOI22D0BWP7T $T=669080 202040 0 0 $X=668790 $Y=201805
X980 89 301 67 298 295 4 3 AOI22D0BWP7T $T=671880 170680 0 0 $X=671590 $Y=170445
X981 95 94 93 67 82 4 3 AOI22D0BWP7T $T=687560 241240 0 180 $X=683910 $Y=237030
X982 88 313 67 290 307 4 3 AOI22D0BWP7T $T=688120 217720 0 0 $X=687830 $Y=217485
X983 88 96 67 97 317 4 3 AOI22D0BWP7T $T=689240 241240 1 0 $X=688950 $Y=237030
X984 90 316 67 307 315 4 3 AOI22D0BWP7T $T=691480 202040 0 0 $X=691190 $Y=201805
X985 86 319 67 315 323 4 3 AOI22D0BWP7T $T=693160 186360 1 0 $X=692870 $Y=182150
X986 89 312 67 323 326 4 3 AOI22D0BWP7T $T=702680 178520 1 0 $X=702390 $Y=174310
X987 86 325 67 327 330 4 3 AOI22D0BWP7T $T=705480 194200 1 0 $X=705190 $Y=189990
X988 90 322 67 317 327 4 3 AOI22D0BWP7T $T=710520 217720 1 180 $X=706870 $Y=217485
X989 86 328 67 331 333 4 3 AOI22D0BWP7T $T=707160 225560 1 0 $X=706870 $Y=221350
X990 85 321 67 326 334 4 3 AOI22D0BWP7T $T=708280 178520 1 0 $X=707990 $Y=174310
X991 90 332 67 103 331 4 3 AOI22D0BWP7T $T=709960 225560 0 0 $X=709670 $Y=225325
X992 89 335 67 330 337 4 3 AOI22D0BWP7T $T=715000 170680 0 0 $X=714710 $Y=170445
X993 85 341 67 343 344 4 3 AOI22D0BWP7T $T=723960 194200 1 0 $X=723670 $Y=189990
X994 89 347 67 333 343 4 3 AOI22D0BWP7T $T=732360 217720 0 0 $X=732070 $Y=217485
X995 85 351 67 337 342 4 3 AOI22D0BWP7T $T=735160 170680 1 0 $X=734870 $Y=166470
X996 85 348 67 108 109 4 3 AOI22D0BWP7T $T=735160 241240 1 0 $X=734870 $Y=237030
X997 3 4 ICV_37 $T=487640 209880 0 0 $X=487350 $Y=209645
X998 3 4 ICV_37 $T=529640 178520 0 0 $X=529350 $Y=178285
X999 3 4 ICV_37 $T=546440 178520 1 0 $X=546150 $Y=174310
X1000 3 4 ICV_37 $T=555400 209880 1 0 $X=555110 $Y=205670
X1001 3 4 ICV_37 $T=571640 170680 0 0 $X=571350 $Y=170445
X1002 3 4 ICV_37 $T=571640 194200 0 0 $X=571350 $Y=193965
X1003 3 4 ICV_37 $T=576120 225560 0 0 $X=575830 $Y=225325
X1004 3 4 ICV_37 $T=595160 170680 0 0 $X=594870 $Y=170445
X1005 3 4 ICV_37 $T=597960 186360 1 0 $X=597670 $Y=182150
X1006 3 4 ICV_37 $T=618120 170680 1 0 $X=617830 $Y=166470
X1007 3 4 ICV_37 $T=627080 209880 0 0 $X=626790 $Y=209645
X1008 3 4 ICV_37 $T=643880 186360 1 0 $X=643590 $Y=182150
X1009 3 4 ICV_37 $T=655640 217720 1 0 $X=655350 $Y=213510
X1010 3 4 ICV_37 $T=664040 194200 0 0 $X=663750 $Y=193965
X1011 3 4 ICV_37 $T=697640 194200 0 0 $X=697350 $Y=193965
X1012 3 4 ICV_37 $T=697640 225560 0 0 $X=697350 $Y=225325
X1013 3 4 ICV_37 $T=702120 194200 1 0 $X=701830 $Y=189990
X1014 3 4 ICV_60 $T=450120 194200 1 0 $X=449830 $Y=189990
X1015 3 4 ICV_60 $T=459080 225560 0 0 $X=458790 $Y=225325
X1016 3 4 ICV_60 $T=478120 186360 0 0 $X=477830 $Y=186125
X1017 3 4 ICV_60 $T=501080 194200 1 0 $X=500790 $Y=189990
X1018 3 4 ICV_60 $T=512280 233400 0 0 $X=511990 $Y=233165
X1019 3 4 ICV_60 $T=512840 186360 1 0 $X=512550 $Y=182150
X1020 3 4 ICV_60 $T=516760 194200 1 0 $X=516470 $Y=189990
X1021 3 4 ICV_60 $T=534120 233400 1 0 $X=533830 $Y=229190
X1022 3 4 ICV_60 $T=576120 194200 0 0 $X=575830 $Y=193965
X1023 3 4 ICV_60 $T=585080 241240 1 0 $X=584790 $Y=237030
X1024 3 4 ICV_60 $T=618120 194200 1 0 $X=617830 $Y=189990
X1025 3 4 ICV_60 $T=618120 217720 1 0 $X=617830 $Y=213510
X1026 3 4 ICV_60 $T=684200 209880 1 0 $X=683910 $Y=205670
X1027 3 4 ICV_60 $T=687000 233400 1 0 $X=686710 $Y=229190
X1028 3 4 ICV_60 $T=687560 170680 1 0 $X=687270 $Y=166470
X1029 3 4 ICV_60 $T=702120 225560 1 0 $X=701830 $Y=221350
X1030 3 4 ICV_60 $T=711080 241240 1 0 $X=710790 $Y=237030
X1031 3 4 ICV_43 $T=450120 186360 1 0 $X=449830 $Y=182150
X1032 3 4 ICV_43 $T=475320 241240 1 0 $X=475030 $Y=237030
X1033 3 4 ICV_43 $T=492120 186360 1 0 $X=491830 $Y=182150
X1034 3 4 ICV_43 $T=492120 217720 0 0 $X=491830 $Y=217485
X1035 3 4 ICV_43 $T=511160 170680 1 0 $X=510870 $Y=166470
X1036 3 4 ICV_43 $T=512280 225560 1 0 $X=511990 $Y=221350
X1037 3 4 ICV_43 $T=534120 209880 0 0 $X=533830 $Y=209645
X1038 3 4 ICV_43 $T=543080 186360 0 0 $X=542790 $Y=186125
X1039 3 4 ICV_43 $T=583960 233400 1 0 $X=583670 $Y=229190
X1040 3 4 ICV_43 $T=594040 162840 0 0 $X=593750 $Y=162605
X1041 3 4 ICV_43 $T=597960 202040 1 0 $X=597670 $Y=197830
X1042 3 4 ICV_43 $T=627080 225560 0 0 $X=626790 $Y=225325
X1043 3 4 ICV_43 $T=648360 186360 0 0 $X=648070 $Y=186125
X1044 3 4 ICV_43 $T=660120 209880 1 0 $X=659830 $Y=205670
X1045 3 4 ICV_43 $T=664600 162840 1 0 $X=664310 $Y=158630
X1046 3 4 ICV_43 $T=688680 202040 0 0 $X=688390 $Y=201805
X1047 3 4 ICV_43 $T=711080 186360 0 0 $X=710790 $Y=186125
X1048 3 4 ICV_43 $T=716120 186360 1 0 $X=715830 $Y=182150
X1049 3 4 ICV_43 $T=717800 209880 0 0 $X=717510 $Y=209645
X1050 3 4 ICV_52 $T=453480 241240 1 0 $X=453190 $Y=237030
X1051 3 4 ICV_52 $T=455720 186360 1 0 $X=455430 $Y=182150
X1052 3 4 ICV_52 $T=459080 178520 1 0 $X=458790 $Y=174310
X1053 3 4 ICV_52 $T=460760 241240 1 0 $X=460470 $Y=237030
X1054 3 4 ICV_52 $T=478680 217720 1 0 $X=478390 $Y=213510
X1055 3 4 ICV_52 $T=487080 170680 0 0 $X=486790 $Y=170445
X1056 3 4 ICV_52 $T=501080 233400 1 0 $X=500790 $Y=229190
X1057 3 4 ICV_52 $T=505560 186360 1 0 $X=505270 $Y=182150
X1058 3 4 ICV_52 $T=534120 178520 1 0 $X=533830 $Y=174310
X1059 3 4 ICV_52 $T=618120 186360 1 0 $X=617830 $Y=182150
X1060 3 4 ICV_52 $T=622040 225560 1 0 $X=621750 $Y=221350
X1061 3 4 ICV_52 $T=645000 217720 0 0 $X=644710 $Y=217485
X1062 3 4 ICV_52 $T=660120 233400 0 0 $X=659830 $Y=233165
X1063 3 4 ICV_52 $T=678040 178520 1 0 $X=677750 $Y=174310
X1064 3 4 ICV_52 $T=697080 186360 0 0 $X=696790 $Y=186125
X1065 3 4 ICV_52 $T=711080 170680 0 0 $X=710790 $Y=170445
X1066 51 3 4 50 BUFFD3BWP7T $T=553720 178520 0 180 $X=549510 $Y=174310
X1067 104 3 4 57 BUFFD3BWP7T $T=722280 202040 0 180 $X=718070 $Y=197830
X1068 105 3 4 99 BUFFD3BWP7T $T=723400 217720 1 180 $X=719190 $Y=217485
X1069 38 118 35 3 4 ND2D1P5BWP7T $T=486520 225560 1 180 $X=482310 $Y=225325
X1070 3 4 ICV_69 $T=449000 178520 1 0 $X=448710 $Y=174310
X1071 3 4 ICV_69 $T=449000 202040 1 0 $X=448710 $Y=197830
X1072 3 4 ICV_69 $T=449000 217720 1 0 $X=448710 $Y=213510
X1073 3 4 ICV_69 $T=449000 225560 0 0 $X=448710 $Y=225325
X1074 3 4 ICV_69 $T=491000 233400 1 0 $X=490710 $Y=229190
X1075 3 4 ICV_69 $T=533000 217720 1 0 $X=532710 $Y=213510
X1076 3 4 ICV_69 $T=575000 170680 0 0 $X=574710 $Y=170445
X1077 3 4 ICV_69 $T=575000 186360 1 0 $X=574710 $Y=182150
X1078 3 4 ICV_69 $T=575000 202040 1 0 $X=574710 $Y=197830
X1079 3 4 ICV_69 $T=575000 209880 1 0 $X=574710 $Y=205670
X1080 3 4 ICV_69 $T=575000 217720 1 0 $X=574710 $Y=213510
X1081 3 4 ICV_69 $T=575000 241240 1 0 $X=574710 $Y=237030
X1082 3 4 ICV_69 $T=617000 209880 0 0 $X=616710 $Y=209645
X1083 3 4 ICV_69 $T=617000 225560 0 0 $X=616710 $Y=225325
X1084 3 4 ICV_69 $T=617000 233400 1 0 $X=616710 $Y=229190
X1085 3 4 ICV_69 $T=659000 217720 1 0 $X=658710 $Y=213510
X1086 3 4 ICV_69 $T=701000 186360 0 0 $X=700710 $Y=186125
X1087 3 4 ICV_69 $T=701000 241240 1 0 $X=700710 $Y=237030
X1088 3 4 17 143 31 ICV_68 $T=485960 178520 0 180 $X=475030 $Y=174310
X1089 3 4 17 144 134 ICV_68 $T=486520 162840 0 180 $X=475590 $Y=158630
X1090 3 4 17 145 32 ICV_68 $T=486520 202040 0 180 $X=475590 $Y=197830
X1091 3 4 45 181 173 ICV_68 $T=527960 233400 1 180 $X=517030 $Y=233165
X1092 3 4 45 179 160 ICV_68 $T=528520 162840 0 180 $X=517590 $Y=158630
X1093 3 4 45 183 174 ICV_68 $T=528520 202040 0 180 $X=517590 $Y=197830
X1094 3 4 45 182 175 ICV_68 $T=528520 209880 1 180 $X=517590 $Y=209645
X1095 3 4 45 192 198 ICV_68 $T=570520 178520 1 180 $X=559590 $Y=178285
X1096 3 4 45 230 238 ICV_68 $T=611400 202040 0 180 $X=600470 $Y=197830
X1097 3 4 45 242 70 ICV_68 $T=611400 225560 1 180 $X=600470 $Y=225325
X1098 3 4 45 229 66 ICV_68 $T=612520 241240 0 180 $X=601590 $Y=237030
X1099 3 4 81 308 297 ICV_68 $T=696520 162840 0 180 $X=685590 $Y=158630
X1100 3 4 81 340 103 ICV_68 $T=726760 241240 0 180 $X=715830 $Y=237030
X1101 3 4 81 339 342 ICV_68 $T=738520 162840 0 180 $X=727590 $Y=158630
X1102 3 4 81 338 337 ICV_68 $T=738520 178520 0 180 $X=727590 $Y=174310
X1103 3 4 81 349 344 ICV_68 $T=738520 186360 1 180 $X=727590 $Y=186125
X1104 3 4 81 350 343 ICV_68 $T=738520 202040 1 180 $X=727590 $Y=201805
X1125 35 49 180 3 4 INR2XD2BWP7T $T=540840 241240 1 0 $X=540550 $Y=237030
.ENDS
***************************************
.SUBCKT ICV_66 1 2
** N=2 EP=2 IP=4 FDC=30
*.SEEDPROM
X0 1 2 DCAP8BWP7T $T=17920 0 0 0 $X=17630 $Y=-235
X1 2 1 DCAP32BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_65 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=26
*.SEEDPROM
X0 2 1 DCAPBWP7T $T=0 0 0 0 $X=-290 $Y=-235
X1 3 4 1 2 5 DFQD0BWP7T $T=12320 0 1 180 $X=1390 $Y=-235
.ENDS
***************************************
.SUBCKT BUFFD4BWP7T I Z VSS VDD
** N=5 EP=4 IP=0 FDC=12
*.SEEDPROM
M0 5 I VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=2080 $Y=345 $D=0
M3 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=2800 $Y=345 $D=0
M4 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=3520 $Y=345 $D=0
M5 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=4240 $Y=345 $D=0
M6 5 I VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M7 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M8 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2080 $Y=2205 $D=16
M9 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=2800 $Y=2205 $D=16
M10 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3520 $Y=2205 $D=16
M11 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=4240 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_51 1 2
** N=2 EP=2 IP=4 FDC=2
*.SEEDPROM
X1 2 1 DCAPBWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT OAI21D2BWP7T B VSS ZN A1 A2 VDD
** N=9 EP=6 IP=0 FDC=12
*.SEEDPROM
M0 VSS B 7 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 7 B VSS VSS N L=1.8e-07 W=1e-06 $X=1345 $Y=345 $D=0
M2 ZN A2 7 VSS N L=1.8e-07 W=1e-06 $X=2080 $Y=345 $D=0
M3 7 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=2800 $Y=345 $D=0
M4 ZN A1 7 VSS N L=1.8e-07 W=1e-06 $X=3520 $Y=345 $D=0
M5 7 A2 ZN VSS N L=1.8e-07 W=1e-06 $X=4240 $Y=345 $D=0
M6 ZN B VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M7 VDD B ZN VDD P L=1.8e-07 W=1.37e-06 $X=1345 $Y=2205 $D=16
M8 8 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2145 $Y=2205 $D=16
M9 ZN A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=2800 $Y=2205 $D=16
M10 9 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3520 $Y=2205 $D=16
M11 VDD A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=4200 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR3D3BWP7T A3 VDD A2 A1 VSS ZN
** N=8 EP=6 IP=0 FDC=30
*.SEEDPROM
M0 ZN A3 VSS VSS N L=1.8e-07 W=6e-07 $X=780 $Y=345 $D=0
M1 VSS A3 ZN VSS N L=1.8e-07 W=6e-07 $X=1500 $Y=345 $D=0
M2 ZN A3 VSS VSS N L=1.8e-07 W=6e-07 $X=2220 $Y=345 $D=0
M3 VSS A3 ZN VSS N L=1.8e-07 W=6e-07 $X=2940 $Y=345 $D=0
M4 ZN A3 VSS VSS N L=1.8e-07 W=6e-07 $X=3660 $Y=345 $D=0
M5 VSS A2 ZN VSS N L=1.8e-07 W=6e-07 $X=4380 $Y=345 $D=0
M6 ZN A2 VSS VSS N L=1.8e-07 W=6e-07 $X=5100 $Y=345 $D=0
M7 VSS A2 ZN VSS N L=1.8e-07 W=6e-07 $X=5820 $Y=345 $D=0
M8 ZN A2 VSS VSS N L=1.8e-07 W=6e-07 $X=6540 $Y=345 $D=0
M9 VSS A2 ZN VSS N L=1.8e-07 W=6e-07 $X=7260 $Y=345 $D=0
M10 ZN A1 VSS VSS N L=1.8e-07 W=6e-07 $X=7980 $Y=345 $D=0
M11 VSS A1 ZN VSS N L=1.8e-07 W=6e-07 $X=8700 $Y=345 $D=0
M12 ZN A1 VSS VSS N L=1.8e-07 W=6e-07 $X=9420 $Y=345 $D=0
M13 VSS A1 ZN VSS N L=1.8e-07 W=6e-07 $X=10140 $Y=345 $D=0
M14 ZN A1 VSS VSS N L=1.8e-07 W=6e-07 $X=10860 $Y=345 $D=0
M15 7 A3 VDD VDD P L=1.8e-07 W=1.36e-06 $X=780 $Y=2215 $D=16
M16 VDD A3 7 VDD P L=1.8e-07 W=1.715e-06 $X=1500 $Y=1860 $D=16
M17 7 A3 VDD VDD P L=1.8e-07 W=1.715e-06 $X=2220 $Y=1860 $D=16
M18 VDD A3 7 VDD P L=1.8e-07 W=1.715e-06 $X=2940 $Y=1860 $D=16
M19 7 A3 VDD VDD P L=1.8e-07 W=1.715e-06 $X=3660 $Y=1860 $D=16
M20 8 A2 7 VDD P L=1.8e-07 W=1.645e-06 $X=4380 $Y=1930 $D=16
M21 7 A2 8 VDD P L=1.8e-07 W=1.645e-06 $X=5100 $Y=1930 $D=16
M22 8 A2 7 VDD P L=1.8e-07 W=1.645e-06 $X=5820 $Y=1930 $D=16
M23 7 A2 8 VDD P L=1.8e-07 W=1.645e-06 $X=6540 $Y=1930 $D=16
M24 8 A2 7 VDD P L=1.8e-07 W=1.645e-06 $X=7260 $Y=1930 $D=16
M25 ZN A1 8 VDD P L=1.8e-07 W=1.715e-06 $X=7980 $Y=1860 $D=16
M26 8 A1 ZN VDD P L=1.8e-07 W=1.715e-06 $X=8700 $Y=1860 $D=16
M27 ZN A1 8 VDD P L=1.8e-07 W=1.715e-06 $X=9420 $Y=1860 $D=16
M28 8 A1 ZN VDD P L=1.8e-07 W=1.715e-06 $X=10140 $Y=1860 $D=16
M29 ZN A1 8 VDD P L=1.8e-07 W=1.36e-06 $X=10860 $Y=2215 $D=16
.ENDS
***************************************
.SUBCKT OR4D1BWP7T A4 A3 A2 A1 VDD VSS Z
** N=11 EP=7 IP=0 FDC=10
*.SEEDPROM
M0 8 A4 VSS VSS N L=1.8e-07 W=5e-07 $X=675 $Y=345 $D=0
M1 VSS A3 8 VSS N L=1.8e-07 W=5e-07 $X=1395 $Y=345 $D=0
M2 8 A2 VSS VSS N L=1.8e-07 W=5e-07 $X=2125 $Y=345 $D=0
M3 VSS A1 8 VSS N L=1.8e-07 W=5e-07 $X=2845 $Y=345 $D=0
M4 Z 8 VSS VSS N L=1.8e-07 W=1e-06 $X=3645 $Y=345 $D=0
M5 9 A4 8 VDD P L=1.8e-07 W=1.37e-06 $X=725 $Y=2205 $D=16
M6 10 A3 9 VDD P L=1.8e-07 W=1.37e-06 $X=1325 $Y=2205 $D=16
M7 11 A2 10 VDD P L=1.8e-07 W=1.37e-06 $X=1925 $Y=2205 $D=16
M8 VDD A1 11 VDD P L=1.8e-07 W=1.37e-06 $X=2525 $Y=2205 $D=16
M9 Z 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3275 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IND3D0BWP7T A1 VSS B1 B2 VDD ZN
** N=9 EP=6 IP=0 FDC=8
*.SEEDPROM
M0 VSS A1 7 VSS N L=1.8e-07 W=4.2e-07 $X=620 $Y=460 $D=0
M1 8 7 VSS VSS N L=1.8e-07 W=5e-07 $X=1340 $Y=460 $D=0
M2 9 B1 8 VSS N L=1.8e-07 W=5e-07 $X=1940 $Y=460 $D=0
M3 ZN B2 9 VSS N L=1.8e-07 W=5e-07 $X=2540 $Y=460 $D=0
M4 VDD A1 7 VDD P L=1.8e-07 W=4.2e-07 $X=620 $Y=2890 $D=16
M5 ZN 7 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1225 $Y=2320 $D=16
M6 VDD B1 ZN VDD P L=1.8e-07 W=6.85e-07 $X=1945 $Y=2320 $D=16
M7 ZN B2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2320 $D=16
.ENDS
***************************************
.SUBCKT IAO21D2BWP7T A1 A2 B ZN VDD VSS
** N=10 EP=6 IP=0 FDC=12
*.SEEDPROM
M0 7 A1 VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS A2 7 VSS N L=1.8e-07 W=1e-06 $X=1345 $Y=345 $D=0
M2 ZN 7 VSS VSS N L=1.8e-07 W=1e-06 $X=2065 $Y=345 $D=0
M3 VSS B ZN VSS N L=1.8e-07 W=1e-06 $X=2785 $Y=345 $D=0
M4 ZN B VSS VSS N L=1.8e-07 W=1e-06 $X=3505 $Y=345 $D=0
M5 VSS 7 ZN VSS N L=1.8e-07 W=1e-06 $X=4225 $Y=345 $D=0
M6 8 A1 7 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M7 VDD A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=1225 $Y=2205 $D=16
M8 9 7 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2125 $Y=2205 $D=16
M9 ZN B 9 VDD P L=1.8e-07 W=1.37e-06 $X=2785 $Y=2205 $D=16
M10 10 B ZN VDD P L=1.8e-07 W=1.37e-06 $X=3505 $Y=2205 $D=16
M11 VDD 7 10 VDD P L=1.8e-07 W=1.37e-06 $X=4225 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OA31D0BWP7T A1 A2 A3 B VSS VDD Z
** N=11 EP=7 IP=0 FDC=10
*.SEEDPROM
M0 8 A1 9 VSS N L=1.8e-07 W=5e-07 $X=665 $Y=750 $D=0
M1 9 A2 8 VSS N L=1.8e-07 W=5e-07 $X=1385 $Y=750 $D=0
M2 8 A3 9 VSS N L=1.8e-07 W=5e-07 $X=2165 $Y=750 $D=0
M3 VSS B 8 VSS N L=1.8e-07 W=5e-07 $X=2910 $Y=750 $D=0
M4 Z 9 VSS VSS N L=1.8e-07 W=5e-07 $X=3670 $Y=750 $D=0
M5 10 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=665 $Y=2860 $D=16
M6 11 A2 10 VDD P L=1.8e-07 W=6.85e-07 $X=1385 $Y=2860 $D=16
M7 9 A3 11 VDD P L=1.8e-07 W=6.85e-07 $X=2105 $Y=2860 $D=16
M8 VDD B 9 VDD P L=1.8e-07 W=6.85e-07 $X=2910 $Y=2860 $D=16
M9 Z 9 VDD VDD P L=1.8e-07 W=6.85e-07 $X=3670 $Y=2860 $D=16
.ENDS
***************************************
.SUBCKT ICV_67 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203
** N=495 EP=201 IP=4556 FDC=10984
*.SEEDPROM
M0 318 335 4 4 N L=1.8e-07 W=1e-06 $X=581240 $Y=357495 $D=0
M1 4 335 318 4 N L=1.8e-07 W=1e-06 $X=581960 $Y=357495 $D=0
M2 318 335 4 4 N L=1.8e-07 W=1e-06 $X=582680 $Y=357495 $D=0
M3 4 102 318 4 N L=1.8e-07 W=1e-06 $X=583400 $Y=357495 $D=0
M4 318 102 4 4 N L=1.8e-07 W=1e-06 $X=584120 $Y=357495 $D=0
M5 4 102 318 4 N L=1.8e-07 W=1e-06 $X=584840 $Y=357495 $D=0
M6 135 107 4 4 N L=1.8e-07 W=5.7e-07 $X=590955 $Y=357925 $D=0
M7 4 107 135 4 N L=1.8e-07 W=5.7e-07 $X=591675 $Y=357925 $D=0
M8 135 107 4 4 N L=1.8e-07 W=5.7e-07 $X=592395 $Y=357925 $D=0
M9 4 107 135 4 N L=1.8e-07 W=5.7e-07 $X=593115 $Y=357925 $D=0
M10 135 107 4 4 N L=1.8e-07 W=5.7e-07 $X=593835 $Y=357925 $D=0
M11 4 107 135 4 N L=1.8e-07 W=5.7e-07 $X=594555 $Y=357925 $D=0
M12 135 107 4 4 N L=1.8e-07 W=5.7e-07 $X=595275 $Y=357925 $D=0
M13 4 101 135 4 N L=1.8e-07 W=5.7e-07 $X=595995 $Y=357925 $D=0
M14 135 101 4 4 N L=1.8e-07 W=5.7e-07 $X=596715 $Y=357925 $D=0
M15 4 101 135 4 N L=1.8e-07 W=5.7e-07 $X=597435 $Y=357925 $D=0
M16 135 101 4 4 N L=1.8e-07 W=5.7e-07 $X=598155 $Y=357925 $D=0
M17 4 101 135 4 N L=1.8e-07 W=5.7e-07 $X=598875 $Y=357925 $D=0
M18 135 101 4 4 N L=1.8e-07 W=5.7e-07 $X=599595 $Y=357925 $D=0
M19 4 101 135 4 N L=1.8e-07 W=5.7e-07 $X=600315 $Y=357925 $D=0
M20 135 102 4 4 N L=1.8e-07 W=5.7e-07 $X=601035 $Y=357925 $D=0
M21 4 102 135 4 N L=1.8e-07 W=5.7e-07 $X=601755 $Y=357925 $D=0
M22 135 102 4 4 N L=1.8e-07 W=5.7e-07 $X=602475 $Y=357925 $D=0
M23 4 102 135 4 N L=1.8e-07 W=5.7e-07 $X=603195 $Y=357925 $D=0
M24 135 102 4 4 N L=1.8e-07 W=5.7e-07 $X=603915 $Y=357925 $D=0
M25 4 102 135 4 N L=1.8e-07 W=5.7e-07 $X=604635 $Y=357925 $D=0
M26 135 102 4 4 N L=1.8e-07 W=5.7e-07 $X=605355 $Y=357925 $D=0
M27 4 134 135 4 N L=1.8e-07 W=5.7e-07 $X=606075 $Y=357925 $D=0
M28 135 134 4 4 N L=1.8e-07 W=5.7e-07 $X=606795 $Y=357925 $D=0
M29 4 134 135 4 N L=1.8e-07 W=5.7e-07 $X=607515 $Y=357925 $D=0
M30 135 134 4 4 N L=1.8e-07 W=5.7e-07 $X=608235 $Y=357925 $D=0
M31 4 134 135 4 N L=1.8e-07 W=5.7e-07 $X=608955 $Y=357925 $D=0
M32 135 134 4 4 N L=1.8e-07 W=5.7e-07 $X=609675 $Y=357925 $D=0
M33 4 134 135 4 N L=1.8e-07 W=5.7e-07 $X=610400 $Y=357925 $D=0
M34 338 335 5 5 P L=1.8e-07 W=1.37e-06 $X=581240 $Y=355265 $D=16
M35 5 335 338 5 P L=1.8e-07 W=1.37e-06 $X=581960 $Y=355265 $D=16
M36 338 335 5 5 P L=1.8e-07 W=1.37e-06 $X=582680 $Y=355265 $D=16
M37 318 102 338 5 P L=1.8e-07 W=1.37e-06 $X=583400 $Y=355265 $D=16
M38 338 102 318 5 P L=1.8e-07 W=1.37e-06 $X=584120 $Y=355265 $D=16
M39 318 102 338 5 P L=1.8e-07 W=1.37e-06 $X=584840 $Y=355265 $D=16
M40 351 107 135 5 P L=1.8e-07 W=1.36e-06 $X=590955 $Y=355265 $D=16
M41 135 107 351 5 P L=1.8e-07 W=1.6e-06 $X=591675 $Y=355265 $D=16
M42 351 107 135 5 P L=1.8e-07 W=1.6e-06 $X=592395 $Y=355265 $D=16
M43 135 107 351 5 P L=1.8e-07 W=1.6e-06 $X=593115 $Y=355265 $D=16
M44 351 107 135 5 P L=1.8e-07 W=1.6e-06 $X=593835 $Y=355265 $D=16
M45 135 107 351 5 P L=1.8e-07 W=1.6e-06 $X=594555 $Y=355265 $D=16
M46 351 107 135 5 P L=1.8e-07 W=1.6e-06 $X=595275 $Y=355265 $D=16
M47 356 101 351 5 P L=1.8e-07 W=1.6e-06 $X=595995 $Y=355265 $D=16
M48 351 101 356 5 P L=1.8e-07 W=1.6e-06 $X=596715 $Y=355265 $D=16
M49 356 101 351 5 P L=1.8e-07 W=1.6e-06 $X=597435 $Y=355265 $D=16
M50 351 101 356 5 P L=1.8e-07 W=1.6e-06 $X=598155 $Y=355265 $D=16
M51 356 101 351 5 P L=1.8e-07 W=1.6e-06 $X=598875 $Y=355265 $D=16
M52 351 101 356 5 P L=1.8e-07 W=1.6e-06 $X=599595 $Y=355265 $D=16
M53 356 101 351 5 P L=1.8e-07 W=1.6e-06 $X=600315 $Y=355265 $D=16
M54 369 102 356 5 P L=1.8e-07 W=1.6e-06 $X=601035 $Y=355265 $D=16
M55 356 102 369 5 P L=1.8e-07 W=1.6e-06 $X=601755 $Y=355265 $D=16
M56 369 102 356 5 P L=1.8e-07 W=1.6e-06 $X=602475 $Y=355265 $D=16
M57 356 102 369 5 P L=1.8e-07 W=1.6e-06 $X=603195 $Y=355265 $D=16
M58 369 102 356 5 P L=1.8e-07 W=1.6e-06 $X=603915 $Y=355265 $D=16
M59 356 102 369 5 P L=1.8e-07 W=1.6e-06 $X=604635 $Y=355265 $D=16
M60 369 102 356 5 P L=1.8e-07 W=1.6e-06 $X=605355 $Y=355265 $D=16
M61 5 134 369 5 P L=1.8e-07 W=1.6e-06 $X=606075 $Y=355265 $D=16
M62 369 134 5 5 P L=1.8e-07 W=1.6e-06 $X=606795 $Y=355265 $D=16
M63 5 134 369 5 P L=1.8e-07 W=1.6e-06 $X=607515 $Y=355265 $D=16
M64 369 134 5 5 P L=1.8e-07 W=1.6e-06 $X=608235 $Y=355265 $D=16
M65 5 134 369 5 P L=1.8e-07 W=1.6e-06 $X=608955 $Y=355265 $D=16
M66 369 134 5 5 P L=1.8e-07 W=1.6e-06 $X=609675 $Y=355265 $D=16
M67 5 134 369 5 P L=1.8e-07 W=1.36e-06 $X=610400 $Y=355265 $D=16
X238 5 4 DCAPBWP7T $T=469160 241240 0 0 $X=468870 $Y=241005
X239 5 4 DCAPBWP7T $T=474760 303960 1 0 $X=474470 $Y=299750
X240 5 4 DCAPBWP7T $T=475320 358840 1 0 $X=475030 $Y=354630
X241 5 4 DCAPBWP7T $T=479240 249080 1 0 $X=478950 $Y=244870
X242 5 4 DCAPBWP7T $T=479240 288280 1 0 $X=478950 $Y=284070
X243 5 4 DCAPBWP7T $T=482040 256920 1 0 $X=481750 $Y=252710
X244 5 4 DCAPBWP7T $T=492120 264760 0 0 $X=491830 $Y=264525
X245 5 4 DCAPBWP7T $T=492120 303960 0 0 $X=491830 $Y=303725
X246 5 4 DCAPBWP7T $T=498840 335320 1 0 $X=498550 $Y=331110
X247 5 4 DCAPBWP7T $T=502760 264760 1 0 $X=502470 $Y=260550
X248 5 4 DCAPBWP7T $T=508360 343160 1 0 $X=508070 $Y=338950
X249 5 4 DCAPBWP7T $T=508920 335320 1 0 $X=508630 $Y=331110
X250 5 4 DCAPBWP7T $T=534120 319640 0 0 $X=533830 $Y=319405
X251 5 4 DCAPBWP7T $T=545880 288280 0 0 $X=545590 $Y=288045
X252 5 4 DCAPBWP7T $T=547560 311800 1 0 $X=547270 $Y=307590
X253 5 4 DCAPBWP7T $T=589560 296120 1 0 $X=589270 $Y=291910
X254 5 4 DCAPBWP7T $T=594040 343160 0 0 $X=593750 $Y=342925
X255 5 4 DCAPBWP7T $T=596280 335320 1 0 $X=595990 $Y=331110
X256 5 4 DCAPBWP7T $T=607480 264760 1 0 $X=607190 $Y=260550
X257 5 4 DCAPBWP7T $T=618120 249080 1 0 $X=617830 $Y=244870
X258 5 4 DCAPBWP7T $T=626520 319640 1 0 $X=626230 $Y=315430
X259 5 4 DCAPBWP7T $T=637720 249080 0 0 $X=637430 $Y=248845
X260 5 4 DCAPBWP7T $T=639400 264760 1 0 $X=639110 $Y=260550
X261 5 4 DCAPBWP7T $T=641080 358840 1 0 $X=640790 $Y=354630
X262 5 4 DCAPBWP7T $T=646120 351000 0 0 $X=645830 $Y=350765
X263 5 4 DCAPBWP7T $T=647800 296120 0 0 $X=647510 $Y=295885
X264 5 4 DCAPBWP7T $T=648920 327480 1 0 $X=648630 $Y=323270
X265 5 4 DCAPBWP7T $T=660120 272600 0 0 $X=659830 $Y=272365
X266 5 4 DCAPBWP7T $T=660120 311800 0 0 $X=659830 $Y=311565
X267 5 4 DCAPBWP7T $T=664040 303960 1 0 $X=663750 $Y=299750
X268 5 4 DCAPBWP7T $T=664600 264760 0 0 $X=664310 $Y=264525
X269 5 4 DCAPBWP7T $T=666840 288280 1 0 $X=666550 $Y=284070
X270 5 4 DCAPBWP7T $T=669080 303960 1 0 $X=668790 $Y=299750
X271 5 4 DCAPBWP7T $T=672440 288280 0 0 $X=672150 $Y=288045
X272 5 4 DCAPBWP7T $T=680280 288280 1 0 $X=679990 $Y=284070
X273 5 4 DCAPBWP7T $T=682520 280440 0 0 $X=682230 $Y=280205
X274 5 4 DCAPBWP7T $T=689800 311800 0 0 $X=689510 $Y=311565
X275 5 4 DCAPBWP7T $T=692600 358840 1 0 $X=692310 $Y=354630
X276 5 4 DCAPBWP7T $T=702120 335320 1 0 $X=701830 $Y=331110
X277 5 4 DCAPBWP7T $T=708840 272600 1 0 $X=708550 $Y=268390
X278 5 4 DCAPBWP7T $T=708840 296120 1 0 $X=708550 $Y=291910
X279 5 4 DCAPBWP7T $T=720040 280440 0 0 $X=719750 $Y=280205
X280 5 4 DCAPBWP7T $T=741320 241240 0 0 $X=741030 $Y=241005
X281 5 4 DCAPBWP7T $T=741320 272600 1 0 $X=741030 $Y=268390
X282 5 4 DCAPBWP7T $T=741320 303960 0 0 $X=741030 $Y=303725
X283 5 4 DCAPBWP7T $T=741320 311800 1 0 $X=741030 $Y=307590
X284 4 5 DCAP8BWP7T $T=450120 256920 1 0 $X=449830 $Y=252710
X285 4 5 DCAP8BWP7T $T=450120 288280 1 0 $X=449830 $Y=284070
X286 4 5 DCAP8BWP7T $T=465800 272600 0 0 $X=465510 $Y=272365
X287 4 5 DCAP8BWP7T $T=469160 303960 0 0 $X=468870 $Y=303725
X288 4 5 DCAP8BWP7T $T=477560 256920 1 0 $X=477270 $Y=252710
X289 4 5 DCAP8BWP7T $T=484840 288280 0 0 $X=484550 $Y=288045
X290 4 5 DCAP8BWP7T $T=485400 319640 1 0 $X=485110 $Y=315430
X291 4 5 DCAP8BWP7T $T=492120 256920 0 0 $X=491830 $Y=256685
X292 4 5 DCAP8BWP7T $T=492120 343160 1 0 $X=491830 $Y=338950
X293 4 5 DCAP8BWP7T $T=495480 303960 1 0 $X=495190 $Y=299750
X294 4 5 DCAP8BWP7T $T=503320 303960 1 0 $X=503030 $Y=299750
X295 4 5 DCAP8BWP7T $T=504440 335320 1 0 $X=504150 $Y=331110
X296 4 5 DCAP8BWP7T $T=510600 280440 1 0 $X=510310 $Y=276230
X297 4 5 DCAP8BWP7T $T=512840 343160 0 0 $X=512550 $Y=342925
X298 4 5 DCAP8BWP7T $T=514520 335320 1 0 $X=514230 $Y=331110
X299 4 5 DCAP8BWP7T $T=515080 264760 0 0 $X=514790 $Y=264525
X300 4 5 DCAP8BWP7T $T=520680 264760 1 0 $X=520390 $Y=260550
X301 4 5 DCAP8BWP7T $T=526840 343160 0 0 $X=526550 $Y=342925
X302 4 5 DCAP8BWP7T $T=527400 256920 1 0 $X=527110 $Y=252710
X303 4 5 DCAP8BWP7T $T=534120 319640 1 0 $X=533830 $Y=315430
X304 4 5 DCAP8BWP7T $T=540840 249080 1 0 $X=540550 $Y=244870
X305 4 5 DCAP8BWP7T $T=541400 358840 1 0 $X=541110 $Y=354630
X306 4 5 DCAP8BWP7T $T=568840 256920 1 0 $X=568550 $Y=252710
X307 4 5 DCAP8BWP7T $T=568840 311800 1 0 $X=568550 $Y=307590
X308 4 5 DCAP8BWP7T $T=576120 249080 1 0 $X=575830 $Y=244870
X309 4 5 DCAP8BWP7T $T=576120 327480 1 0 $X=575830 $Y=323270
X310 4 5 DCAP8BWP7T $T=576120 358840 1 0 $X=575830 $Y=354630
X311 4 5 DCAP8BWP7T $T=583960 288280 1 0 $X=583670 $Y=284070
X312 4 5 DCAP8BWP7T $T=585640 358840 1 0 $X=585350 $Y=354630
X313 4 5 DCAP8BWP7T $T=591240 264760 1 0 $X=590950 $Y=260550
X314 4 5 DCAP8BWP7T $T=610840 335320 1 0 $X=610550 $Y=331110
X315 4 5 DCAP8BWP7T $T=610840 343160 0 0 $X=610550 $Y=342925
X316 4 5 DCAP8BWP7T $T=611400 319640 0 0 $X=611110 $Y=319405
X317 4 5 DCAP8BWP7T $T=611400 358840 1 0 $X=611110 $Y=354630
X318 4 5 DCAP8BWP7T $T=618120 303960 1 0 $X=617830 $Y=299750
X319 4 5 DCAP8BWP7T $T=618120 311800 0 0 $X=617830 $Y=311565
X320 4 5 DCAP8BWP7T $T=618120 327480 0 0 $X=617830 $Y=327245
X321 4 5 DCAP8BWP7T $T=618120 343160 0 0 $X=617830 $Y=342925
X322 4 5 DCAP8BWP7T $T=621480 272600 0 0 $X=621190 $Y=272365
X323 4 5 DCAP8BWP7T $T=622040 319640 1 0 $X=621750 $Y=315430
X324 4 5 DCAP8BWP7T $T=622600 358840 1 0 $X=622310 $Y=354630
X325 4 5 DCAP8BWP7T $T=623720 272600 1 0 $X=623430 $Y=268390
X326 4 5 DCAP8BWP7T $T=631000 311800 1 0 $X=630710 $Y=307590
X327 4 5 DCAP8BWP7T $T=634920 264760 1 0 $X=634630 $Y=260550
X328 4 5 DCAP8BWP7T $T=653400 296120 0 0 $X=653110 $Y=295885
X329 4 5 DCAP8BWP7T $T=653400 327480 1 0 $X=653110 $Y=323270
X330 4 5 DCAP8BWP7T $T=654520 288280 0 0 $X=654230 $Y=288045
X331 4 5 DCAP8BWP7T $T=660120 264760 0 0 $X=659830 $Y=264525
X332 4 5 DCAP8BWP7T $T=664040 272600 0 0 $X=663750 $Y=272365
X333 4 5 DCAP8BWP7T $T=666280 249080 0 0 $X=665990 $Y=248845
X334 4 5 DCAP8BWP7T $T=685320 311800 0 0 $X=685030 $Y=311565
X335 4 5 DCAP8BWP7T $T=694840 351000 0 0 $X=694550 $Y=350765
X336 4 5 DCAP8BWP7T $T=702120 241240 0 0 $X=701830 $Y=241005
X337 4 5 DCAP8BWP7T $T=702120 327480 1 0 $X=701830 $Y=323270
X338 4 5 DCAP8BWP7T $T=712200 343160 1 0 $X=711910 $Y=338950
X339 4 5 DCAP8BWP7T $T=715000 351000 0 0 $X=714710 $Y=350765
X340 4 5 DCAP8BWP7T $T=737400 280440 0 0 $X=737110 $Y=280205
X341 4 5 DCAP8BWP7T $T=737400 343160 0 0 $X=737110 $Y=342925
X342 4 5 DCAP8BWP7T $T=738520 264760 0 0 $X=738230 $Y=264525
X343 4 5 DCAP8BWP7T $T=738520 272600 0 0 $X=738230 $Y=272365
X344 4 5 DCAP8BWP7T $T=738520 288280 0 0 $X=738230 $Y=288045
X345 4 5 DCAP8BWP7T $T=738520 296120 0 0 $X=738230 $Y=295885
X346 4 5 DCAP8BWP7T $T=738520 311800 0 0 $X=738230 $Y=311565
X347 4 5 DCAP8BWP7T $T=738520 319640 1 0 $X=738230 $Y=315430
X348 4 5 DCAP8BWP7T $T=738520 327480 1 0 $X=738230 $Y=323270
X349 4 5 DCAP8BWP7T $T=738520 343160 1 0 $X=738230 $Y=338950
X350 4 5 DCAP8BWP7T $T=738520 351000 1 0 $X=738230 $Y=346790
X351 4 5 DCAP8BWP7T $T=738520 358840 1 0 $X=738230 $Y=354630
X352 4 5 DCAP4BWP7T $T=450120 256920 0 0 $X=449830 $Y=256685
X353 4 5 DCAP4BWP7T $T=450120 343160 0 0 $X=449830 $Y=342925
X354 4 5 DCAP4BWP7T $T=488200 351000 0 0 $X=487910 $Y=350765
X355 4 5 DCAP4BWP7T $T=488760 358840 1 0 $X=488470 $Y=354630
X356 4 5 DCAP4BWP7T $T=534120 327480 0 0 $X=533830 $Y=327245
X357 4 5 DCAP4BWP7T $T=534120 351000 1 0 $X=533830 $Y=346790
X358 4 5 DCAP4BWP7T $T=546440 319640 1 0 $X=546150 $Y=315430
X359 4 5 DCAP4BWP7T $T=572760 311800 0 0 $X=572470 $Y=311565
X360 4 5 DCAP4BWP7T $T=576120 311800 1 0 $X=575830 $Y=307590
X361 4 5 DCAP4BWP7T $T=614200 241240 0 0 $X=613910 $Y=241005
X362 4 5 DCAP4BWP7T $T=614200 256920 1 0 $X=613910 $Y=252710
X363 4 5 DCAP4BWP7T $T=614200 264760 0 0 $X=613910 $Y=264525
X364 4 5 DCAP4BWP7T $T=614200 280440 1 0 $X=613910 $Y=276230
X365 4 5 DCAP4BWP7T $T=614760 303960 0 0 $X=614470 $Y=303725
X366 4 5 DCAP4BWP7T $T=618120 256920 1 0 $X=617830 $Y=252710
X367 4 5 DCAP4BWP7T $T=618120 272600 1 0 $X=617830 $Y=268390
X368 4 5 DCAP4BWP7T $T=656200 303960 1 0 $X=655910 $Y=299750
X369 4 5 DCAP4BWP7T $T=660120 249080 0 0 $X=659830 $Y=248845
X370 4 5 DCAP4BWP7T $T=678600 319640 1 0 $X=678310 $Y=315430
X371 4 5 DCAP4BWP7T $T=687000 249080 1 0 $X=686710 $Y=244870
X372 4 5 DCAP4BWP7T $T=702120 249080 0 0 $X=701830 $Y=248845
X373 4 5 DCAP4BWP7T $T=702120 311800 0 0 $X=701830 $Y=311565
X374 4 5 DCAP4BWP7T $T=702120 343160 0 0 $X=701830 $Y=342925
X375 4 5 DCAP4BWP7T $T=702120 351000 0 0 $X=701830 $Y=350765
X376 4 5 DCAP4BWP7T $T=711080 351000 1 0 $X=710790 $Y=346790
X377 4 5 DCAP4BWP7T $T=729560 303960 1 0 $X=729270 $Y=299750
X378 4 5 DCAP4BWP7T $T=740200 296120 1 0 $X=739910 $Y=291910
X379 4 5 DCAP4BWP7T $T=740760 335320 0 0 $X=740470 $Y=335085
X380 4 5 ICV_40 $T=450120 241240 0 0 $X=449830 $Y=241005
X381 4 5 ICV_40 $T=450120 249080 1 0 $X=449830 $Y=244870
X382 4 5 ICV_40 $T=450120 311800 1 0 $X=449830 $Y=307590
X383 4 5 ICV_40 $T=450120 343160 1 0 $X=449830 $Y=338950
X384 4 5 ICV_40 $T=459080 256920 1 0 $X=458790 $Y=252710
X385 4 5 ICV_40 $T=459080 264760 0 0 $X=458790 $Y=264525
X386 4 5 ICV_40 $T=460200 288280 1 0 $X=459910 $Y=284070
X387 4 5 ICV_40 $T=468040 303960 1 0 $X=467750 $Y=299750
X388 4 5 ICV_40 $T=468040 327480 0 0 $X=467750 $Y=327245
X389 4 5 ICV_40 $T=471400 249080 0 0 $X=471110 $Y=248845
X390 4 5 ICV_40 $T=482600 241240 0 0 $X=482310 $Y=241005
X391 4 5 ICV_40 $T=482600 296120 1 0 $X=482310 $Y=291910
X392 4 5 ICV_40 $T=483160 280440 1 0 $X=482870 $Y=276230
X393 4 5 ICV_40 $T=483160 343160 0 0 $X=482870 $Y=342925
X394 4 5 ICV_40 $T=483720 264760 0 0 $X=483430 $Y=264525
X395 4 5 ICV_40 $T=483720 288280 1 0 $X=483430 $Y=284070
X396 4 5 ICV_40 $T=483720 296120 0 0 $X=483430 $Y=295885
X397 4 5 ICV_40 $T=484280 249080 1 0 $X=483990 $Y=244870
X398 4 5 ICV_40 $T=484280 335320 1 0 $X=483990 $Y=331110
X399 4 5 ICV_40 $T=492120 272600 1 0 $X=491830 $Y=268390
X400 4 5 ICV_40 $T=492120 288280 0 0 $X=491830 $Y=288045
X401 4 5 ICV_40 $T=492120 335320 1 0 $X=491830 $Y=331110
X402 4 5 ICV_40 $T=492120 351000 0 0 $X=491830 $Y=350765
X403 4 5 ICV_40 $T=496040 264760 1 0 $X=495750 $Y=260550
X404 4 5 ICV_40 $T=501640 343160 1 0 $X=501350 $Y=338950
X405 4 5 ICV_40 $T=515080 303960 0 0 $X=514790 $Y=303725
X406 4 5 ICV_40 $T=524600 241240 0 0 $X=524310 $Y=241005
X407 4 5 ICV_40 $T=524600 311800 0 0 $X=524310 $Y=311565
X408 4 5 ICV_40 $T=525720 335320 1 0 $X=525430 $Y=331110
X409 4 5 ICV_40 $T=526280 358840 1 0 $X=525990 $Y=354630
X410 4 5 ICV_40 $T=534120 327480 1 0 $X=533830 $Y=323270
X411 4 5 ICV_40 $T=539160 288280 1 0 $X=538870 $Y=284070
X412 4 5 ICV_40 $T=539160 288280 0 0 $X=538870 $Y=288045
X413 4 5 ICV_40 $T=548680 335320 1 0 $X=548390 $Y=331110
X414 4 5 ICV_40 $T=552040 272600 1 0 $X=551750 $Y=268390
X415 4 5 ICV_40 $T=553160 249080 1 0 $X=552870 $Y=244870
X416 4 5 ICV_40 $T=555400 303960 1 0 $X=555110 $Y=299750
X417 4 5 ICV_40 $T=567160 241240 0 0 $X=566870 $Y=241005
X418 4 5 ICV_40 $T=567160 264760 0 0 $X=566870 $Y=264525
X419 4 5 ICV_40 $T=567160 272600 0 0 $X=566870 $Y=272365
X420 4 5 ICV_40 $T=567160 319640 1 0 $X=566870 $Y=315430
X421 4 5 ICV_40 $T=567720 296120 1 0 $X=567430 $Y=291910
X422 4 5 ICV_40 $T=567720 351000 1 0 $X=567430 $Y=346790
X423 4 5 ICV_40 $T=568280 280440 1 0 $X=567990 $Y=276230
X424 4 5 ICV_40 $T=576120 272600 0 0 $X=575830 $Y=272365
X425 4 5 ICV_40 $T=576120 311800 0 0 $X=575830 $Y=311565
X426 4 5 ICV_40 $T=576120 335320 0 0 $X=575830 $Y=335085
X427 4 5 ICV_40 $T=579480 264760 1 0 $X=579190 $Y=260550
X428 4 5 ICV_40 $T=585080 249080 0 0 $X=584790 $Y=248845
X429 4 5 ICV_40 $T=589560 335320 1 0 $X=589270 $Y=331110
X430 4 5 ICV_40 $T=608600 288280 0 0 $X=608310 $Y=288045
X431 4 5 ICV_40 $T=609160 327480 0 0 $X=608870 $Y=327245
X432 4 5 ICV_40 $T=618120 343160 1 0 $X=617830 $Y=338950
X433 4 5 ICV_40 $T=618120 351000 0 0 $X=617830 $Y=350765
X434 4 5 ICV_40 $T=627080 335320 0 0 $X=626790 $Y=335085
X435 4 5 ICV_40 $T=634360 358840 1 0 $X=634070 $Y=354630
X436 4 5 ICV_40 $T=636040 256920 0 0 $X=635750 $Y=256685
X437 4 5 ICV_40 $T=641080 296120 0 0 $X=640790 $Y=295885
X438 4 5 ICV_40 $T=650600 249080 1 0 $X=650310 $Y=244870
X439 4 5 ICV_40 $T=651720 319640 1 0 $X=651430 $Y=315430
X440 4 5 ICV_40 $T=651720 335320 1 0 $X=651430 $Y=331110
X441 4 5 ICV_40 $T=652280 256920 0 0 $X=651990 $Y=256685
X442 4 5 ICV_40 $T=652280 288280 1 0 $X=651990 $Y=284070
X443 4 5 ICV_40 $T=660120 288280 1 0 $X=659830 $Y=284070
X444 4 5 ICV_40 $T=660120 327480 1 0 $X=659830 $Y=323270
X445 4 5 ICV_40 $T=669640 264760 0 0 $X=669350 $Y=264525
X446 4 5 ICV_40 $T=671320 327480 1 0 $X=671030 $Y=323270
X447 4 5 ICV_40 $T=672440 272600 0 0 $X=672150 $Y=272365
X448 4 5 ICV_40 $T=678040 311800 1 0 $X=677750 $Y=307590
X449 4 5 ICV_40 $T=684760 288280 1 0 $X=684470 $Y=284070
X450 4 5 ICV_40 $T=685880 358840 1 0 $X=685590 $Y=354630
X451 4 5 ICV_40 $T=687000 296120 1 0 $X=686710 $Y=291910
X452 4 5 ICV_40 $T=692600 264760 1 0 $X=692310 $Y=260550
X453 4 5 ICV_40 $T=692600 319640 1 0 $X=692310 $Y=315430
X454 4 5 ICV_40 $T=693160 256920 1 0 $X=692870 $Y=252710
X455 4 5 ICV_40 $T=693720 311800 0 0 $X=693430 $Y=311565
X456 4 5 ICV_40 $T=694280 343160 1 0 $X=693990 $Y=338950
X457 4 5 ICV_40 $T=702120 272600 1 0 $X=701830 $Y=268390
X458 4 5 ICV_40 $T=702120 296120 1 0 $X=701830 $Y=291910
X459 4 5 ICV_40 $T=702120 335320 0 0 $X=701830 $Y=335085
X460 4 5 ICV_40 $T=711080 311800 1 0 $X=710790 $Y=307590
X461 4 5 ICV_40 $T=711080 319640 0 0 $X=710790 $Y=319405
X462 4 5 ICV_40 $T=720600 343160 1 0 $X=720310 $Y=338950
X463 4 5 ICV_40 $T=727880 288280 0 0 $X=727590 $Y=288045
X464 4 5 ICV_40 $T=734600 303960 0 0 $X=734310 $Y=303725
X465 4 5 ICV_40 $T=735160 249080 1 0 $X=734870 $Y=244870
X466 4 5 ICV_40 $T=735160 256920 1 0 $X=734870 $Y=252710
X467 4 5 ICV_40 $T=735160 264760 1 0 $X=734870 $Y=260550
X468 4 5 ICV_40 $T=735720 256920 0 0 $X=735430 $Y=256685
X469 4 5 ICV_40 $T=735720 303960 1 0 $X=735430 $Y=299750
X470 5 4 DCAP64BWP7T $T=450120 280440 0 0 $X=449830 $Y=280205
X471 5 4 DCAP64BWP7T $T=450120 311800 0 0 $X=449830 $Y=311565
X472 5 4 DCAP64BWP7T $T=492120 311800 1 0 $X=491830 $Y=307590
X473 5 4 DCAP64BWP7T $T=492120 351000 1 0 $X=491830 $Y=346790
X474 5 4 DCAP64BWP7T $T=534120 351000 0 0 $X=533830 $Y=350765
X475 5 4 DCAP64BWP7T $T=576120 351000 0 0 $X=575830 $Y=350765
X476 5 4 DCAP64BWP7T $T=618120 280440 0 0 $X=617830 $Y=280205
X477 5 4 DCAP64BWP7T $T=618120 303960 0 0 $X=617830 $Y=303725
X478 5 4 DCAP64BWP7T $T=660120 303960 0 0 $X=659830 $Y=303725
X479 5 4 DCAP64BWP7T $T=660120 319640 0 0 $X=659830 $Y=319405
X480 5 4 DCAP64BWP7T $T=702120 327480 0 0 $X=701830 $Y=327245
X522 5 4 DCAP32BWP7T $T=450120 249080 0 0 $X=449830 $Y=248845
X523 5 4 DCAP32BWP7T $T=450120 303960 1 0 $X=449830 $Y=299750
X524 5 4 DCAP32BWP7T $T=450120 327480 0 0 $X=449830 $Y=327245
X525 5 4 DCAP32BWP7T $T=450120 335320 0 0 $X=449830 $Y=335085
X526 5 4 DCAP32BWP7T $T=465800 296120 0 0 $X=465510 $Y=295885
X527 5 4 DCAP32BWP7T $T=492120 272600 0 0 $X=491830 $Y=272365
X528 5 4 DCAP32BWP7T $T=492120 311800 0 0 $X=491830 $Y=311565
X529 5 4 DCAP32BWP7T $T=534120 272600 1 0 $X=533830 $Y=268390
X530 5 4 DCAP32BWP7T $T=543640 264760 1 0 $X=543350 $Y=260550
X531 5 4 DCAP32BWP7T $T=550360 280440 1 0 $X=550070 $Y=276230
X532 5 4 DCAP32BWP7T $T=576120 343160 1 0 $X=575830 $Y=338950
X533 5 4 DCAP32BWP7T $T=576120 343160 0 0 $X=575830 $Y=342925
X534 5 4 DCAP32BWP7T $T=581720 288280 0 0 $X=581430 $Y=288045
X535 5 4 DCAP32BWP7T $T=594600 296120 1 0 $X=594310 $Y=291910
X536 5 4 DCAP32BWP7T $T=595160 288280 1 0 $X=594870 $Y=284070
X537 5 4 DCAP32BWP7T $T=596280 264760 0 0 $X=595990 $Y=264525
X538 5 4 DCAP32BWP7T $T=618120 256920 0 0 $X=617830 $Y=256685
X539 5 4 DCAP32BWP7T $T=618120 264760 0 0 $X=617830 $Y=264525
X540 5 4 DCAP32BWP7T $T=625960 343160 0 0 $X=625670 $Y=342925
X541 5 4 DCAP32BWP7T $T=660120 241240 0 0 $X=659830 $Y=241005
X542 5 4 DCAP32BWP7T $T=660120 311800 1 0 $X=659830 $Y=307590
X543 5 4 DCAP32BWP7T $T=662920 343160 0 0 $X=662630 $Y=342925
X544 5 4 DCAP32BWP7T $T=674680 264760 1 0 $X=674390 $Y=260550
X545 5 4 DCAP32BWP7T $T=676360 343160 1 0 $X=676070 $Y=338950
X546 5 4 DCAP32BWP7T $T=681400 249080 0 0 $X=681110 $Y=248845
X547 5 4 DCAP32BWP7T $T=683080 351000 1 0 $X=682790 $Y=346790
X548 5 4 DCAP32BWP7T $T=702120 256920 1 0 $X=701830 $Y=252710
X549 5 4 DCAP32BWP7T $T=702120 264760 0 0 $X=701830 $Y=264525
X550 5 4 DCAP32BWP7T $T=702120 280440 0 0 $X=701830 $Y=280205
X551 5 4 DCAP32BWP7T $T=702120 303960 0 0 $X=701830 $Y=303725
X552 5 4 DCAP32BWP7T $T=702120 358840 1 0 $X=701830 $Y=354630
X553 5 4 DCAP32BWP7T $T=709960 241240 0 0 $X=709670 $Y=241005
X554 5 4 DCAP32BWP7T $T=711640 319640 1 0 $X=711350 $Y=315430
X555 5 4 DCAP32BWP7T $T=716680 351000 1 0 $X=716390 $Y=346790
X556 5 4 DCAP32BWP7T $T=723400 311800 1 0 $X=723110 $Y=307590
X557 393 4 5 385 INVD1BWP7T $T=642760 358840 1 0 $X=642470 $Y=354630
X558 291 4 5 78 CKBD0BWP7T $T=539160 288280 1 180 $X=536630 $Y=288045
X684 277 4 44 66 5 ND2D1BWP7T $T=516200 319640 0 0 $X=515910 $Y=319405
X685 277 4 67 69 5 ND2D1BWP7T $T=518440 319640 0 0 $X=518150 $Y=319405
X686 76 4 75 73 5 ND2D1BWP7T $T=528520 249080 0 180 $X=525990 $Y=244870
X687 288 4 38 73 5 ND2D1BWP7T $T=528520 264760 0 180 $X=525990 $Y=260550
X688 288 4 35 74 5 ND2D1BWP7T $T=528520 280440 0 180 $X=525990 $Y=276230
X689 277 4 63 74 5 ND2D1BWP7T $T=526280 319640 0 0 $X=525990 $Y=319405
X690 277 4 55 73 5 ND2D1BWP7T $T=528520 327480 0 180 $X=525990 $Y=323270
X691 288 4 48 77 5 ND2D1BWP7T $T=537480 280440 1 180 $X=534950 $Y=280205
X692 277 4 34 77 5 ND2D1BWP7T $T=538040 319640 1 180 $X=535510 $Y=319405
X693 288 4 40 82 5 ND2D1BWP7T $T=536920 288280 1 0 $X=536630 $Y=284070
X694 277 4 36 82 5 ND2D1BWP7T $T=541960 319640 0 180 $X=539430 $Y=315430
X695 277 4 72 84 5 ND2D1BWP7T $T=541960 327480 1 0 $X=541670 $Y=323270
X696 288 4 65 85 5 ND2D1BWP7T $T=542520 249080 0 0 $X=542230 $Y=248845
X697 288 4 31 66 5 ND2D1BWP7T $T=546440 303960 0 180 $X=543910 $Y=299750
X698 277 4 47 85 5 ND2D1BWP7T $T=544200 327480 1 0 $X=543910 $Y=323270
X699 76 4 87 85 5 ND2D1BWP7T $T=545320 249080 1 0 $X=545030 $Y=244870
X700 288 4 49 69 5 ND2D1BWP7T $T=549800 288280 1 180 $X=547270 $Y=288045
X701 288 4 15 84 5 ND2D1BWP7T $T=550920 319640 0 180 $X=548390 $Y=315430
X702 76 4 96 74 5 ND2D1BWP7T $T=553160 249080 0 180 $X=550630 $Y=244870
X703 66 4 105 318 5 ND2D1BWP7T $T=563240 303960 1 0 $X=562950 $Y=299750
X704 69 4 108 318 5 ND2D1BWP7T $T=576680 303960 0 0 $X=576390 $Y=303725
X705 74 4 112 318 5 ND2D1BWP7T $T=576680 319640 0 0 $X=576390 $Y=319405
X706 77 4 99 318 5 ND2D1BWP7T $T=581160 319640 1 180 $X=578630 $Y=319405
X707 73 4 111 318 5 ND2D1BWP7T $T=581720 327480 1 0 $X=581430 $Y=323270
X708 82 4 130 318 5 ND2D1BWP7T $T=603560 319640 1 0 $X=603270 $Y=315430
X709 318 4 365 84 5 ND2D1BWP7T $T=628200 319640 0 0 $X=627910 $Y=319405
X710 85 4 154 318 5 ND2D1BWP7T $T=646680 311800 0 180 $X=644150 $Y=307590
X711 135 4 170 84 5 ND2D1BWP7T $T=654520 241240 1 180 $X=651990 $Y=241005
X712 135 4 165 85 5 ND2D1BWP7T $T=652280 264760 1 0 $X=651990 $Y=260550
X713 135 4 411 77 5 ND2D1BWP7T $T=652280 311800 0 0 $X=651990 $Y=311565
X714 160 4 173 84 5 ND2D1BWP7T $T=660680 351000 0 0 $X=660390 $Y=350765
X715 135 4 176 74 5 ND2D1BWP7T $T=661800 272600 0 0 $X=661510 $Y=272365
X716 135 4 178 73 5 ND2D1BWP7T $T=678600 327480 1 0 $X=678310 $Y=323270
X717 160 4 185 74 5 ND2D1BWP7T $T=683080 351000 0 180 $X=680550 $Y=346790
X718 160 4 188 73 5 ND2D1BWP7T $T=685880 358840 0 180 $X=683350 $Y=354630
X719 160 4 179 77 5 ND2D1BWP7T $T=691480 351000 1 180 $X=688950 $Y=350765
X720 135 4 423 69 5 ND2D1BWP7T $T=693720 311800 1 180 $X=691190 $Y=311565
X721 160 4 193 85 5 ND2D1BWP7T $T=692600 351000 0 0 $X=692310 $Y=350765
X722 160 4 195 66 5 ND2D1BWP7T $T=694280 358840 1 0 $X=693990 $Y=354630
X746 110 4 5 300 INVD0BWP7T $T=578360 335320 0 180 $X=576390 $Y=331110
X747 36 210 11 209 4 5 OAI21D0BWP7T $T=455160 343160 1 180 $X=452070 $Y=342925
X748 10 218 15 216 4 5 OAI21D0BWP7T $T=452920 303960 0 0 $X=452630 $Y=303725
X749 10 220 31 219 4 5 OAI21D0BWP7T $T=465800 296120 1 180 $X=462710 $Y=295885
X750 10 215 35 212 4 5 OAI21D0BWP7T $T=471400 249080 1 180 $X=468310 $Y=248845
X751 10 39 38 211 4 5 OAI21D0BWP7T $T=473640 241240 1 180 $X=470550 $Y=241005
X752 37 226 40 233 4 5 OAI21D0BWP7T $T=470840 272600 0 0 $X=470550 $Y=272365
X753 47 46 11 229 4 5 OAI21D0BWP7T $T=479800 358840 0 180 $X=476710 $Y=354630
X754 37 230 35 236 4 5 OAI21D0BWP7T $T=478120 249080 0 0 $X=477830 $Y=248845
X755 37 225 48 234 4 5 OAI21D0BWP7T $T=479240 264760 1 0 $X=478950 $Y=260550
X756 37 237 49 235 4 5 OAI21D0BWP7T $T=483720 288280 0 180 $X=480630 $Y=284070
X757 35 52 50 245 4 5 OAI21D0BWP7T $T=483720 256920 1 0 $X=483430 $Y=252710
X758 40 248 50 243 4 5 OAI21D0BWP7T $T=495480 280440 0 180 $X=492390 $Y=276230
X759 37 239 31 249 4 5 OAI21D0BWP7T $T=492680 303960 1 0 $X=492390 $Y=299750
X760 38 254 50 259 4 5 OAI21D0BWP7T $T=494920 256920 1 0 $X=494630 $Y=252710
X761 55 256 11 262 4 5 OAI21D0BWP7T $T=498840 343160 1 0 $X=498550 $Y=338950
X762 37 238 15 246 4 5 OAI21D0BWP7T $T=504440 319640 0 0 $X=504150 $Y=319405
X763 48 268 50 255 4 5 OAI21D0BWP7T $T=510600 280440 0 180 $X=507510 $Y=276230
X764 31 270 50 261 4 5 OAI21D0BWP7T $T=508920 303960 1 0 $X=508630 $Y=299750
X765 49 269 50 260 4 5 OAI21D0BWP7T $T=513960 288280 0 180 $X=510870 $Y=284070
X766 63 273 11 286 4 5 OAI21D0BWP7T $T=518440 343160 0 0 $X=518150 $Y=342925
X767 50 278 15 284 4 5 OAI21D0BWP7T $T=524600 311800 1 180 $X=521510 $Y=311565
X768 11 274 72 287 4 5 OAI21D0BWP7T $T=524040 343160 0 0 $X=523750 $Y=342925
X769 89 297 90 92 4 5 OAI21D0BWP7T $T=547000 351000 1 0 $X=546710 $Y=346790
X770 302 304 99 309 4 5 OAI21D0BWP7T $T=555400 272600 0 0 $X=555110 $Y=272365
X771 99 306 320 319 4 5 OAI21D0BWP7T $T=564920 296120 1 0 $X=564630 $Y=291910
X772 106 314 99 323 4 5 OAI21D0BWP7T $T=566040 256920 1 0 $X=565750 $Y=252710
X773 316 301 108 321 4 5 OAI21D0BWP7T $T=568840 311800 0 180 $X=565750 $Y=307590
X774 316 322 99 312 4 5 OAI21D0BWP7T $T=567160 319640 0 0 $X=566870 $Y=319405
X775 302 299 111 332 4 5 OAI21D0BWP7T $T=576680 264760 1 0 $X=576390 $Y=260550
X776 302 311 112 330 4 5 OAI21D0BWP7T $T=576680 280440 0 0 $X=576390 $Y=280205
X777 108 298 320 331 4 5 OAI21D0BWP7T $T=576680 296120 0 0 $X=576390 $Y=295885
X778 111 337 320 327 4 5 OAI21D0BWP7T $T=584520 303960 0 180 $X=581430 $Y=299750
X779 118 313 99 339 4 5 OAI21D0BWP7T $T=582280 256920 0 0 $X=581990 $Y=256685
X780 112 345 320 328 4 5 OAI21D0BWP7T $T=591240 303960 1 180 $X=588150 $Y=303725
X781 316 349 111 347 4 5 OAI21D0BWP7T $T=595720 327480 0 180 $X=592630 $Y=323270
X782 316 346 112 343 4 5 OAI21D0BWP7T $T=600760 335320 0 180 $X=597670 $Y=331110
X783 302 348 108 359 4 5 OAI21D0BWP7T $T=601320 264760 1 0 $X=601030 $Y=260550
X784 302 344 105 360 4 5 OAI21D0BWP7T $T=602440 272600 0 0 $X=602150 $Y=272365
X785 105 355 320 361 4 5 OAI21D0BWP7T $T=603000 303960 0 0 $X=602710 $Y=303725
X786 118 358 365 368 4 5 OAI21D0BWP7T $T=606920 256920 1 0 $X=606630 $Y=252710
X787 316 353 105 371 4 5 OAI21D0BWP7T $T=609720 311800 1 0 $X=609430 $Y=307590
X788 302 357 365 376 4 5 OAI21D0BWP7T $T=618680 272600 0 0 $X=618390 $Y=272365
X789 365 373 320 372 4 5 OAI21D0BWP7T $T=621480 288280 0 180 $X=618390 $Y=284070
X790 316 362 365 379 4 5 OAI21D0BWP7T $T=619240 327480 1 0 $X=618950 $Y=323270
X791 302 384 130 383 4 5 OAI21D0BWP7T $T=625960 272600 0 0 $X=625670 $Y=272365
X792 116 392 365 148 4 5 OAI21D0BWP7T $T=634360 241240 1 180 $X=631270 $Y=241005
X793 316 388 130 387 4 5 OAI21D0BWP7T $T=634360 319640 0 180 $X=631270 $Y=315430
X794 106 390 365 375 4 5 OAI21D0BWP7T $T=634920 256920 0 180 $X=631830 $Y=252710
X795 130 389 320 386 4 5 OAI21D0BWP7T $T=636600 311800 1 0 $X=636310 $Y=307590
X796 302 402 154 397 4 5 OAI21D0BWP7T $T=643880 264760 0 180 $X=640790 $Y=260550
X797 154 404 320 401 4 5 OAI21D0BWP7T $T=646120 296120 0 180 $X=643030 $Y=291910
X798 316 403 154 400 4 5 OAI21D0BWP7T $T=646120 311800 1 180 $X=643030 $Y=311565
X799 156 405 165 407 4 5 OAI21D0BWP7T $T=649480 256920 0 0 $X=649190 $Y=256685
X800 156 412 411 409 4 5 OAI21D0BWP7T $T=654520 288280 1 180 $X=651430 $Y=288045
X801 156 413 178 419 4 5 OAI21D0BWP7T $T=665720 280440 1 0 $X=665430 $Y=276230
X802 168 416 179 425 4 5 OAI21D0BWP7T $T=666280 351000 0 0 $X=665990 $Y=350765
X803 156 418 423 426 4 5 OAI21D0BWP7T $T=666840 319640 1 0 $X=666550 $Y=315430
X804 411 424 164 432 4 5 OAI21D0BWP7T $T=668520 288280 1 0 $X=668230 $Y=284070
X805 156 427 176 421 4 5 OAI21D0BWP7T $T=669640 272600 0 0 $X=669350 $Y=272365
X806 179 415 184 430 4 5 OAI21D0BWP7T $T=673560 343160 1 0 $X=673270 $Y=338950
X807 156 434 186 187 4 5 OAI21D0BWP7T $T=678600 241240 0 0 $X=678310 $Y=241005
X808 178 435 164 438 4 5 OAI21D0BWP7T $T=679720 272600 0 0 $X=679430 $Y=272365
X809 423 437 164 417 4 5 OAI21D0BWP7T $T=683640 319640 0 180 $X=680550 $Y=315430
X810 175 431 411 440 4 5 OAI21D0BWP7T $T=681960 288280 1 0 $X=681670 $Y=284070
X811 175 442 423 447 4 5 OAI21D0BWP7T $T=687560 288280 0 0 $X=687270 $Y=288045
X812 176 446 164 190 4 5 OAI21D0BWP7T $T=692040 249080 0 180 $X=688950 $Y=244870
X813 171 455 411 451 4 5 OAI21D0BWP7T $T=696520 296120 0 180 $X=693430 $Y=291910
X814 168 448 188 443 4 5 OAI21D0BWP7T $T=705480 343160 0 180 $X=702390 $Y=338950
X815 168 459 185 462 4 5 OAI21D0BWP7T $T=704360 343160 0 0 $X=704070 $Y=342925
X816 186 197 164 450 4 5 OAI21D0BWP7T $T=709960 241240 1 180 $X=706870 $Y=241005
X817 167 465 411 457 4 5 OAI21D0BWP7T $T=711640 319640 0 180 $X=708550 $Y=315430
X818 185 463 184 468 4 5 OAI21D0BWP7T $T=709400 343160 1 0 $X=709110 $Y=338950
X819 171 469 423 464 4 5 OAI21D0BWP7T $T=713320 272600 0 180 $X=710230 $Y=268390
X820 411 461 163 476 4 5 OAI21D0BWP7T $T=710520 296120 1 0 $X=710230 $Y=291910
X821 175 467 178 454 4 5 OAI21D0BWP7T $T=716120 256920 1 180 $X=713030 $Y=256685
X822 171 460 178 473 4 5 OAI21D0BWP7T $T=718920 249080 1 180 $X=715830 $Y=248845
X823 167 482 423 485 4 5 OAI21D0BWP7T $T=722840 303960 0 0 $X=722550 $Y=303725
X824 167 483 178 480 4 5 OAI21D0BWP7T $T=726200 264760 0 180 $X=723110 $Y=260550
X825 168 484 195 479 4 5 OAI21D0BWP7T $T=725080 358840 1 0 $X=724790 $Y=354630
X826 423 492 163 495 4 5 OAI21D0BWP7T $T=734600 280440 0 0 $X=734310 $Y=280205
X827 195 494 184 486 4 5 OAI21D0BWP7T $T=738520 351000 0 180 $X=735430 $Y=346790
X874 4 5 DCAP16BWP7T $T=450120 264760 0 0 $X=449830 $Y=264525
X875 4 5 DCAP16BWP7T $T=450120 296120 1 0 $X=449830 $Y=291910
X876 4 5 DCAP16BWP7T $T=450120 319640 0 0 $X=449830 $Y=319405
X877 4 5 DCAP16BWP7T $T=450120 351000 1 0 $X=449830 $Y=346790
X878 4 5 DCAP16BWP7T $T=461320 343160 1 0 $X=461030 $Y=338950
X879 4 5 DCAP16BWP7T $T=468040 264760 1 0 $X=467750 $Y=260550
X880 4 5 DCAP16BWP7T $T=473640 296120 1 0 $X=473350 $Y=291910
X881 4 5 DCAP16BWP7T $T=475320 335320 1 0 $X=475030 $Y=331110
X882 4 5 DCAP16BWP7T $T=479800 358840 1 0 $X=479510 $Y=354630
X883 4 5 DCAP16BWP7T $T=480360 303960 1 0 $X=480070 $Y=299750
X884 4 5 DCAP16BWP7T $T=481480 272600 1 0 $X=481190 $Y=268390
X885 4 5 DCAP16BWP7T $T=482040 264760 1 0 $X=481750 $Y=260550
X886 4 5 DCAP16BWP7T $T=492120 241240 0 0 $X=491830 $Y=241005
X887 4 5 DCAP16BWP7T $T=492120 319640 0 0 $X=491830 $Y=319405
X888 4 5 DCAP16BWP7T $T=506120 303960 0 0 $X=505830 $Y=303725
X889 4 5 DCAP16BWP7T $T=507240 319640 0 0 $X=506950 $Y=319405
X890 4 5 DCAP16BWP7T $T=515640 241240 0 0 $X=515350 $Y=241005
X891 4 5 DCAP16BWP7T $T=520680 343160 1 0 $X=520390 $Y=338950
X892 4 5 DCAP16BWP7T $T=522360 272600 0 0 $X=522070 $Y=272365
X893 4 5 DCAP16BWP7T $T=523480 264760 0 0 $X=523190 $Y=264525
X894 4 5 DCAP16BWP7T $T=523480 303960 1 0 $X=523190 $Y=299750
X895 4 5 DCAP16BWP7T $T=534120 303960 1 0 $X=533830 $Y=299750
X896 4 5 DCAP16BWP7T $T=534120 335320 0 0 $X=533830 $Y=335085
X897 4 5 DCAP16BWP7T $T=546440 272600 0 0 $X=546150 $Y=272365
X898 4 5 DCAP16BWP7T $T=546440 303960 1 0 $X=546150 $Y=299750
X899 4 5 DCAP16BWP7T $T=549800 288280 0 0 $X=549510 $Y=288045
X900 4 5 DCAP16BWP7T $T=550920 319640 1 0 $X=550630 $Y=315430
X901 4 5 DCAP16BWP7T $T=550920 358840 1 0 $X=550630 $Y=354630
X902 4 5 DCAP16BWP7T $T=556520 256920 1 0 $X=556230 $Y=252710
X903 4 5 DCAP16BWP7T $T=558200 241240 0 0 $X=557910 $Y=241005
X904 4 5 DCAP16BWP7T $T=558200 272600 0 0 $X=557910 $Y=272365
X905 4 5 DCAP16BWP7T $T=562680 249080 0 0 $X=562390 $Y=248845
X906 4 5 DCAP16BWP7T $T=564920 358840 1 0 $X=564630 $Y=354630
X907 4 5 DCAP16BWP7T $T=565480 296120 0 0 $X=565190 $Y=295885
X908 4 5 DCAP16BWP7T $T=565480 303960 1 0 $X=565190 $Y=299750
X909 4 5 DCAP16BWP7T $T=576120 249080 0 0 $X=575830 $Y=248845
X910 4 5 DCAP16BWP7T $T=576120 264760 0 0 $X=575830 $Y=264525
X911 4 5 DCAP16BWP7T $T=576120 280440 1 0 $X=575830 $Y=276230
X912 4 5 DCAP16BWP7T $T=581160 319640 0 0 $X=580870 $Y=319405
X913 4 5 DCAP16BWP7T $T=584520 303960 1 0 $X=584230 $Y=299750
X914 4 5 DCAP16BWP7T $T=591240 303960 0 0 $X=590950 $Y=303725
X915 4 5 DCAP16BWP7T $T=605240 241240 0 0 $X=604950 $Y=241005
X916 4 5 DCAP16BWP7T $T=605800 303960 0 0 $X=605510 $Y=303725
X917 4 5 DCAP16BWP7T $T=608040 319640 1 0 $X=607750 $Y=315430
X918 4 5 DCAP16BWP7T $T=618120 241240 0 0 $X=617830 $Y=241005
X919 4 5 DCAP16BWP7T $T=618120 249080 0 0 $X=617830 $Y=248845
X920 4 5 DCAP16BWP7T $T=618120 280440 1 0 $X=617830 $Y=276230
X921 4 5 DCAP16BWP7T $T=618120 319640 0 0 $X=617830 $Y=319405
X922 4 5 DCAP16BWP7T $T=618120 335320 0 0 $X=617830 $Y=335085
X923 4 5 DCAP16BWP7T $T=628200 343160 1 0 $X=627910 $Y=338950
X924 4 5 DCAP16BWP7T $T=629880 351000 0 0 $X=629590 $Y=350765
X925 4 5 DCAP16BWP7T $T=632120 288280 1 0 $X=631830 $Y=284070
X926 4 5 DCAP16BWP7T $T=633240 272600 1 0 $X=632950 $Y=268390
X927 4 5 DCAP16BWP7T $T=641640 249080 1 0 $X=641350 $Y=244870
X928 4 5 DCAP16BWP7T $T=642760 288280 0 0 $X=642470 $Y=288045
X929 4 5 DCAP16BWP7T $T=642760 335320 1 0 $X=642470 $Y=331110
X930 4 5 DCAP16BWP7T $T=646120 296120 1 0 $X=645830 $Y=291910
X931 4 5 DCAP16BWP7T $T=646680 272600 0 0 $X=646390 $Y=272365
X932 4 5 DCAP16BWP7T $T=646680 311800 1 0 $X=646390 $Y=307590
X933 4 5 DCAP16BWP7T $T=646680 327480 0 0 $X=646390 $Y=327245
X934 4 5 DCAP16BWP7T $T=647240 303960 1 0 $X=646950 $Y=299750
X935 4 5 DCAP16BWP7T $T=648360 319640 0 0 $X=648070 $Y=319405
X936 4 5 DCAP16BWP7T $T=650040 249080 0 0 $X=649750 $Y=248845
X937 4 5 DCAP16BWP7T $T=660120 351000 1 0 $X=659830 $Y=346790
X938 4 5 DCAP16BWP7T $T=679720 280440 1 0 $X=679430 $Y=276230
X939 4 5 DCAP16BWP7T $T=681400 241240 0 0 $X=681110 $Y=241005
X940 4 5 DCAP16BWP7T $T=690360 288280 0 0 $X=690070 $Y=288045
X941 4 5 DCAP16BWP7T $T=690360 343160 0 0 $X=690070 $Y=342925
X942 4 5 DCAP16BWP7T $T=692040 249080 1 0 $X=691750 $Y=244870
X943 4 5 DCAP16BWP7T $T=702120 256920 0 0 $X=701830 $Y=256685
X944 4 5 DCAP16BWP7T $T=702120 311800 1 0 $X=701830 $Y=307590
X945 4 5 DCAP16BWP7T $T=702120 319640 0 0 $X=701830 $Y=319405
X946 4 5 DCAP16BWP7T $T=702120 351000 1 0 $X=701830 $Y=346790
X947 4 5 DCAP16BWP7T $T=714440 264760 1 0 $X=714150 $Y=260550
X948 4 5 DCAP16BWP7T $T=714440 288280 1 0 $X=714150 $Y=284070
X949 4 5 DCAP16BWP7T $T=715560 272600 0 0 $X=715270 $Y=272365
X950 4 5 DCAP16BWP7T $T=716120 256920 0 0 $X=715830 $Y=256685
X951 4 5 DCAP16BWP7T $T=717240 327480 1 0 $X=716950 $Y=323270
X952 4 5 DCAP16BWP7T $T=720600 303960 1 0 $X=720310 $Y=299750
X953 4 5 DCAP16BWP7T $T=725080 280440 0 0 $X=724790 $Y=280205
X954 4 5 DCAP16BWP7T $T=726200 264760 1 0 $X=725910 $Y=260550
X955 4 5 DCAP16BWP7T $T=731240 296120 1 0 $X=730950 $Y=291910
X1005 305 288 5 4 INVD2BWP7T $T=557080 319640 1 180 $X=554550 $Y=319405
X1062 7 210 4 5 6 DFQD0BWP7T $T=461320 351000 1 180 $X=450390 $Y=350765
X1063 7 12 4 5 29 DFQD0BWP7T $T=451240 296120 0 0 $X=450950 $Y=295885
X1064 13 215 4 5 9 DFQD0BWP7T $T=463000 256920 1 180 $X=452070 $Y=256685
X1065 13 17 4 5 20 DFQD0BWP7T $T=452920 272600 1 0 $X=452630 $Y=268390
X1066 7 218 4 5 22 DFQD0BWP7T $T=468040 311800 0 180 $X=457110 $Y=307590
X1067 7 220 4 5 30 DFQD0BWP7T $T=473640 296120 0 180 $X=462710 $Y=291910
X1068 13 230 4 5 222 DFQD0BWP7T $T=477560 256920 0 180 $X=466630 $Y=252710
X1069 13 225 4 5 213 DFQD0BWP7T $T=466920 264760 0 0 $X=466630 $Y=264525
X1070 7 238 4 5 224 DFQD0BWP7T $T=485400 319640 0 180 $X=474470 $Y=315430
X1071 7 241 4 5 42 DFQD0BWP7T $T=486520 327480 1 180 $X=475590 $Y=327245
X1072 58 254 4 5 53 DFQD0BWP7T $T=503320 249080 0 180 $X=492390 $Y=244870
X1073 7 250 4 5 266 DFQD0BWP7T $T=492680 327480 0 0 $X=492390 $Y=327245
X1074 58 248 4 5 240 DFQD0BWP7T $T=506120 280440 1 180 $X=495190 $Y=280205
X1075 7 256 4 5 258 DFQD0BWP7T $T=495480 343160 0 0 $X=495190 $Y=342925
X1076 7 54 4 5 56 DFQD0BWP7T $T=496040 358840 1 0 $X=495750 $Y=354630
X1077 58 268 4 5 242 DFQD0BWP7T $T=509480 272600 0 180 $X=498550 $Y=268390
X1078 58 269 4 5 252 DFQD0BWP7T $T=509480 296120 0 180 $X=498550 $Y=291910
X1079 7 270 4 5 257 DFQD0BWP7T $T=509480 319640 0 180 $X=498550 $Y=315430
X1080 58 64 4 5 61 DFQD0BWP7T $T=515640 241240 1 180 $X=504710 $Y=241005
X1081 7 273 4 5 282 DFQD0BWP7T $T=510040 343160 1 0 $X=509750 $Y=338950
X1082 7 274 4 5 68 DFQD0BWP7T $T=510040 358840 1 0 $X=509750 $Y=354630
X1083 58 278 4 5 253 DFQD0BWP7T $T=521240 311800 1 180 $X=510310 $Y=311565
X1084 58 281 4 5 265 DFQD0BWP7T $T=523480 303960 0 180 $X=512550 $Y=299750
X1085 7 272 4 5 275 DFQD0BWP7T $T=512840 327480 0 0 $X=512550 $Y=327245
X1086 58 279 4 5 276 DFQD0BWP7T $T=527960 249080 1 180 $X=517030 $Y=248845
X1087 58 285 4 5 263 DFQD0BWP7T $T=545880 256920 1 180 $X=534950 $Y=256685
X1088 58 295 4 5 289 DFQD0BWP7T $T=547000 351000 0 180 $X=536070 $Y=346790
X1089 58 293 4 5 290 DFQD0BWP7T $T=550920 296120 1 180 $X=539990 $Y=295885
X1090 58 298 4 5 303 DFQD0BWP7T $T=545880 288280 1 0 $X=545590 $Y=284070
X1091 58 299 4 5 308 DFQD0BWP7T $T=547560 264760 0 0 $X=547270 $Y=264525
X1092 58 306 4 5 310 DFQD0BWP7T $T=554840 296120 0 0 $X=554550 $Y=295885
X1093 58 311 4 5 324 DFQD0BWP7T $T=558760 280440 0 0 $X=558470 $Y=280205
X1094 58 313 4 5 325 DFQD0BWP7T $T=559320 256920 0 0 $X=559030 $Y=256685
X1095 58 304 4 5 317 DFQD0BWP7T $T=559320 272600 1 0 $X=559030 $Y=268390
X1096 58 314 4 5 326 DFQD0BWP7T $T=559880 249080 1 0 $X=559590 $Y=244870
X1097 58 115 4 5 340 DFQD0BWP7T $T=576680 241240 0 0 $X=576390 $Y=241005
X1098 58 345 4 5 334 DFQD0BWP7T $T=593480 311800 1 180 $X=582550 $Y=311565
X1099 58 346 4 5 329 DFQD0BWP7T $T=594040 335320 1 180 $X=583110 $Y=335085
X1100 58 348 4 5 342 DFQD0BWP7T $T=596280 264760 1 180 $X=585350 $Y=264525
X1101 58 344 4 5 352 DFQD0BWP7T $T=586200 280440 1 0 $X=585910 $Y=276230
X1102 58 349 4 5 350 DFQD0BWP7T $T=605800 343160 0 180 $X=594870 $Y=338950
X1103 58 353 4 5 364 DFQD0BWP7T $T=596280 311800 0 0 $X=595990 $Y=311565
X1104 58 355 4 5 363 DFQD0BWP7T $T=596840 303960 1 0 $X=596550 $Y=299750
X1105 58 362 4 5 354 DFQD0BWP7T $T=609160 327480 1 180 $X=598230 $Y=327245
X1106 58 357 4 5 367 DFQD0BWP7T $T=599080 280440 1 0 $X=598790 $Y=276230
X1107 58 358 4 5 370 DFQD0BWP7T $T=600760 249080 0 0 $X=600470 $Y=248845
X1108 149 384 4 5 378 DFQD0BWP7T $T=632120 288280 0 180 $X=621190 $Y=284070
X1109 149 388 4 5 381 DFQD0BWP7T $T=634360 327480 1 180 $X=623430 $Y=327245
X1110 149 390 4 5 380 DFQD0BWP7T $T=634920 264760 0 180 $X=623990 $Y=260550
X1111 149 392 4 5 141 DFQD0BWP7T $T=637720 249080 1 180 $X=626790 $Y=248845
X1112 149 373 4 5 377 DFQD0BWP7T $T=642760 288280 1 180 $X=631830 $Y=288045
X1113 149 403 4 5 394 DFQD0BWP7T $T=646680 327480 1 180 $X=635750 $Y=327245
X1114 149 402 4 5 395 DFQD0BWP7T $T=647240 280440 0 180 $X=636310 $Y=276230
X1115 149 399 4 5 406 DFQD0BWP7T $T=637160 343160 1 0 $X=636870 $Y=338950
X1116 149 415 4 5 429 DFQD0BWP7T $T=662920 343160 1 0 $X=662630 $Y=338950
X1117 149 416 4 5 183 DFQD0BWP7T $T=664040 358840 1 0 $X=663750 $Y=354630
X1118 149 424 4 5 414 DFQD0BWP7T $T=670760 303960 1 0 $X=670470 $Y=299750
X1119 149 431 4 5 436 DFQD0BWP7T $T=674120 288280 0 0 $X=673830 $Y=288045
X1120 149 435 4 5 428 DFQD0BWP7T $T=676360 264760 0 0 $X=676070 $Y=264525
X1121 149 445 4 5 433 DFQD0BWP7T $T=692600 327480 0 180 $X=681670 $Y=323270
X1122 149 446 4 5 180 DFQD0BWP7T $T=693160 256920 0 180 $X=682230 $Y=252710
X1123 149 442 4 5 422 DFQD0BWP7T $T=685880 311800 1 0 $X=685590 $Y=307590
X1124 149 448 4 5 189 DFQD0BWP7T $T=696520 335320 1 180 $X=685590 $Y=335085
X1125 149 460 4 5 449 DFQD0BWP7T $T=704360 249080 0 0 $X=704070 $Y=248845
X1126 149 461 4 5 471 DFQD0BWP7T $T=704360 311800 0 0 $X=704070 $Y=311565
X1127 149 459 4 5 199 DFQD0BWP7T $T=704360 351000 0 0 $X=704070 $Y=350765
X1128 149 469 4 5 452 DFQD0BWP7T $T=715560 272600 1 180 $X=704630 $Y=272365
X1129 149 465 4 5 456 DFQD0BWP7T $T=717240 303960 0 180 $X=706310 $Y=299750
X1130 149 458 4 5 441 DFQD0BWP7T $T=717240 327480 0 180 $X=706310 $Y=323270
X1131 149 483 4 5 474 DFQD0BWP7T $T=727880 272600 0 180 $X=716950 $Y=268390
X1132 149 466 4 5 470 DFQD0BWP7T $T=729000 319640 1 180 $X=718070 $Y=319405
X1133 149 463 4 5 472 DFQD0BWP7T $T=729000 335320 0 180 $X=718070 $Y=331110
X1134 149 203 4 5 200 DFQD0BWP7T $T=735160 249080 0 180 $X=724230 $Y=244870
X1135 149 490 4 5 201 DFQD0BWP7T $T=735720 256920 1 180 $X=724790 $Y=256685
X1136 149 492 4 5 488 DFQD0BWP7T $T=738520 272600 1 180 $X=727590 $Y=272365
X1137 149 491 4 5 489 DFQD0BWP7T $T=738520 296120 1 180 $X=727590 $Y=295885
X1138 149 478 4 5 477 DFQD0BWP7T $T=738520 311800 1 180 $X=727590 $Y=311565
X1139 149 493 4 5 487 DFQD0BWP7T $T=738520 327480 0 180 $X=727590 $Y=323270
X1140 149 494 4 5 481 DFQD0BWP7T $T=738520 343160 0 180 $X=727590 $Y=338950
X1141 149 484 4 5 202 DFQD0BWP7T $T=738520 358840 0 180 $X=727590 $Y=354630
X1142 58 322 4 5 307 DFQD1BWP7T $T=569960 335320 0 180 $X=559030 $Y=331110
X1143 149 405 4 5 152 DFQD1BWP7T $T=650040 249080 1 180 $X=639110 $Y=248845
X1144 149 418 4 5 410 DFQD1BWP7T $T=672440 327480 1 180 $X=661510 $Y=327245
X1145 149 427 4 5 174 DFQD1BWP7T $T=674680 264760 0 180 $X=663750 $Y=260550
X1146 149 434 4 5 181 DFQD1BWP7T $T=681400 249080 1 180 $X=670470 $Y=248845
X1147 86 43 4 5 BUFFD1P5BWP7T $T=547000 343160 0 180 $X=543910 $Y=338950
X1148 297 95 4 5 BUFFD1P5BWP7T $T=553720 319640 1 180 $X=550630 $Y=319405
X1149 307 100 4 5 BUFFD1P5BWP7T $T=556520 335320 1 0 $X=556230 $Y=331110
X1150 142 144 4 5 BUFFD1P5BWP7T $T=622600 311800 0 0 $X=622310 $Y=311565
X1151 410 166 4 5 BUFFD1P5BWP7T $T=653400 327480 0 180 $X=650310 $Y=323270
X1152 292 277 5 4 CKND2BWP7T $T=539720 335320 0 180 $X=537190 $Y=331110
X1153 329 4 5 113 CKBD1BWP7T $T=580600 335320 0 180 $X=578070 $Y=331110
X1154 364 4 5 131 CKBD1BWP7T $T=608040 319640 0 180 $X=605510 $Y=315430
X1155 354 4 5 133 CKBD1BWP7T $T=610840 335320 0 180 $X=608310 $Y=331110
X1156 350 4 5 127 CKBD1BWP7T $T=611960 343160 0 180 $X=609430 $Y=338950
X1157 381 4 5 146 CKBD1BWP7T $T=628200 343160 0 180 $X=625670 $Y=338950
X1158 394 4 5 151 CKBD1BWP7T $T=636040 335320 1 180 $X=633510 $Y=335085
X1159 157 4 5 160 CKBD1BWP7T $T=647800 351000 0 0 $X=647510 $Y=350765
X1160 8 33 5 4 33 214 34 MAOI22D0BWP7T $T=464120 319640 0 0 $X=463830 $Y=319405
X1161 217 33 5 4 33 227 36 MAOI22D0BWP7T $T=470840 319640 1 0 $X=470550 $Y=315430
X1162 28 33 5 4 33 223 44 MAOI22D0BWP7T $T=473640 343160 1 0 $X=473350 $Y=338950
X1163 42 33 5 4 33 241 67 MAOI22D0BWP7T $T=482600 335320 0 0 $X=482310 $Y=335085
X1164 228 33 5 4 33 232 47 MAOI22D0BWP7T $T=482600 351000 1 0 $X=482310 $Y=346790
X1165 266 33 5 4 33 250 55 MAOI22D0BWP7T $T=504440 335320 0 180 $X=500230 $Y=331110
X1166 251 267 5 4 267 271 35 MAOI22D0BWP7T $T=504440 264760 1 0 $X=504150 $Y=260550
X1167 275 33 5 4 33 272 63 MAOI22D0BWP7T $T=514520 335320 0 180 $X=510310 $Y=331110
X1168 276 267 5 4 267 279 65 MAOI22D0BWP7T $T=514520 256920 1 0 $X=514230 $Y=252710
X1169 244 267 5 4 267 280 40 MAOI22D0BWP7T $T=519000 280440 1 0 $X=518710 $Y=276230
X1170 263 267 5 4 267 285 38 MAOI22D0BWP7T $T=519560 264760 0 0 $X=519270 $Y=264525
X1171 264 267 5 4 267 283 49 MAOI22D0BWP7T $T=524040 288280 0 0 $X=523750 $Y=288045
X1172 265 267 5 4 267 281 31 MAOI22D0BWP7T $T=534680 296120 0 0 $X=534390 $Y=295885
X1173 289 33 5 4 33 295 72 MAOI22D0BWP7T $T=534680 343160 1 0 $X=534390 $Y=338950
X1174 290 267 5 4 267 293 15 MAOI22D0BWP7T $T=537480 303960 0 0 $X=537190 $Y=303725
X1175 247 267 5 4 267 294 48 MAOI22D0BWP7T $T=546440 280440 1 0 $X=546150 $Y=276230
X1176 143 125 5 4 125 138 365 MAOI22D0BWP7T $T=623720 249080 0 180 $X=619510 $Y=244870
X1177 433 192 5 4 192 445 179 MAOI22D0BWP7T $T=692600 327480 1 0 $X=692310 $Y=323270
X1178 441 192 5 4 192 458 188 MAOI22D0BWP7T $T=707720 335320 0 180 $X=703510 $Y=331110
X1179 470 192 5 4 192 466 185 MAOI22D0BWP7T $T=713880 335320 1 180 $X=709670 $Y=335085
X1180 477 169 5 4 169 478 411 MAOI22D0BWP7T $T=723400 311800 0 180 $X=719190 $Y=307590
X1181 489 169 5 4 169 491 423 MAOI22D0BWP7T $T=735720 303960 0 180 $X=731510 $Y=299750
X1182 201 169 5 4 169 490 178 MAOI22D0BWP7T $T=738520 264760 1 180 $X=734310 $Y=264525
X1183 487 192 5 4 192 493 195 MAOI22D0BWP7T $T=734600 319640 1 0 $X=734310 $Y=315430
X1184 101 107 366 134 92 4 5 OAI31D1BWP7T $T=606920 343160 0 0 $X=606630 $Y=342925
X1185 137 124 374 139 92 4 5 OAI31D1BWP7T $T=618680 358840 1 0 $X=618390 $Y=354630
X1186 10 14 18 20 221 5 4 AOI22D0BWP7T $T=453480 272600 0 0 $X=453190 $Y=272365
X1187 10 21 18 23 213 5 4 AOI22D0BWP7T $T=455720 256920 1 0 $X=455430 $Y=252710
X1188 10 211 18 25 32 5 4 AOI22D0BWP7T $T=456840 241240 0 0 $X=456550 $Y=241005
X1189 10 212 18 9 222 5 4 AOI22D0BWP7T $T=457960 249080 1 0 $X=457670 $Y=244870
X1190 11 209 26 6 217 5 4 AOI22D0BWP7T $T=457960 343160 1 0 $X=457670 $Y=338950
X1191 10 216 26 22 224 5 4 AOI22D0BWP7T $T=465800 303960 0 0 $X=465510 $Y=303725
X1192 10 219 26 30 231 5 4 AOI22D0BWP7T $T=466920 288280 1 0 $X=466630 $Y=284070
X1193 11 229 26 41 228 5 4 AOI22D0BWP7T $T=471960 358840 1 0 $X=471670 $Y=354630
X1194 37 233 26 221 240 5 4 AOI22D0BWP7T $T=479800 280440 1 0 $X=479510 $Y=276230
X1195 37 234 18 213 242 5 4 AOI22D0BWP7T $T=480360 264760 0 0 $X=480070 $Y=264525
X1196 37 236 18 222 51 5 4 AOI22D0BWP7T $T=480920 249080 1 0 $X=480630 $Y=244870
X1197 50 243 18 240 244 5 4 AOI22D0BWP7T $T=483160 272600 0 0 $X=482870 $Y=272365
X1198 50 245 24 51 251 5 4 AOI22D0BWP7T $T=492680 264760 1 0 $X=492390 $Y=260550
X1199 37 235 26 3 252 5 4 AOI22D0BWP7T $T=492680 296120 1 0 $X=492390 $Y=291910
X1200 37 246 26 224 253 5 4 AOI22D0BWP7T $T=492680 319640 1 0 $X=492390 $Y=315430
X1201 50 255 24 242 247 5 4 AOI22D0BWP7T $T=497160 264760 1 180 $X=493510 $Y=264525
X1202 37 249 26 231 257 5 4 AOI22D0BWP7T $T=493800 303960 0 0 $X=493510 $Y=303725
X1203 50 259 24 53 263 5 4 AOI22D0BWP7T $T=498840 256920 0 0 $X=498550 $Y=256685
X1204 59 57 26 56 258 5 4 AOI22D0BWP7T $T=502200 351000 1 180 $X=498550 $Y=350765
X1205 50 260 26 252 264 5 4 AOI22D0BWP7T $T=499400 288280 0 0 $X=499110 $Y=288045
X1206 50 261 26 257 265 5 4 AOI22D0BWP7T $T=499960 303960 1 0 $X=499670 $Y=299750
X1207 50 62 24 61 276 5 4 AOI22D0BWP7T $T=505560 249080 0 0 $X=505270 $Y=248845
X1208 11 262 26 258 266 5 4 AOI22D0BWP7T $T=512840 343160 1 180 $X=509190 $Y=342925
X1209 11 286 26 282 275 5 4 AOI22D0BWP7T $T=522360 335320 1 0 $X=522070 $Y=331110
X1210 50 284 26 253 290 5 4 AOI22D0BWP7T $T=522920 303960 0 0 $X=522630 $Y=303725
X1211 59 71 26 70 282 5 4 AOI22D0BWP7T $T=526280 358840 0 180 $X=522630 $Y=354630
X1212 11 287 26 68 289 5 4 AOI22D0BWP7T $T=525160 351000 0 0 $X=524870 $Y=350765
X1213 310 312 100 315 316 5 4 AOI22D0BWP7T $T=560440 319640 0 0 $X=560150 $Y=319405
X1214 320 319 317 310 315 5 4 AOI22D0BWP7T $T=566600 288280 1 180 $X=562950 $Y=288045
X1215 303 321 104 315 316 5 4 AOI22D0BWP7T $T=567160 319640 0 180 $X=563510 $Y=315430
X1216 302 309 315 317 325 5 4 AOI22D0BWP7T $T=580040 272600 0 180 $X=576390 $Y=268390
X1217 320 327 308 333 315 5 4 AOI22D0BWP7T $T=578360 288280 0 0 $X=578070 $Y=288045
X1218 320 328 324 334 315 5 4 AOI22D0BWP7T $T=578360 311800 1 0 $X=578070 $Y=307590
X1219 302 332 315 308 114 5 4 AOI22D0BWP7T $T=582280 256920 1 180 $X=578630 $Y=256685
X1220 116 117 24 340 128 5 4 AOI22D0BWP7T $T=581160 249080 1 0 $X=580870 $Y=244870
X1221 302 330 315 324 119 5 4 AOI22D0BWP7T $T=586760 272600 1 180 $X=583110 $Y=272365
X1222 334 343 113 315 316 5 4 AOI22D0BWP7T $T=587320 327480 0 180 $X=583670 $Y=323270
X1223 118 339 315 325 326 5 4 AOI22D0BWP7T $T=591240 264760 0 180 $X=587590 $Y=260550
X1224 333 347 127 315 316 5 4 AOI22D0BWP7T $T=590120 319640 0 0 $X=589830 $Y=319405
X1225 320 331 342 303 315 5 4 AOI22D0BWP7T $T=594600 296120 0 180 $X=590950 $Y=291910
X1226 106 323 315 326 340 5 4 AOI22D0BWP7T $T=596840 264760 1 0 $X=596550 $Y=260550
X1227 302 359 315 342 132 5 4 AOI22D0BWP7T $T=604120 264760 1 0 $X=603830 $Y=260550
X1228 118 368 315 370 380 5 4 AOI22D0BWP7T $T=609160 264760 1 0 $X=608870 $Y=260550
X1229 302 360 315 352 136 5 4 AOI22D0BWP7T $T=609160 272600 0 0 $X=608870 $Y=272365
X1230 320 361 352 363 315 5 4 AOI22D0BWP7T $T=609160 303960 1 0 $X=608870 $Y=299750
X1231 363 371 131 315 316 5 4 AOI22D0BWP7T $T=618680 319640 1 0 $X=618390 $Y=315430
X1232 367 372 377 315 320 5 4 AOI22D0BWP7T $T=619800 296120 0 0 $X=619510 $Y=295885
X1233 106 375 315 380 141 5 4 AOI22D0BWP7T $T=620360 256920 1 0 $X=620070 $Y=252710
X1234 302 376 315 367 370 5 4 AOI22D0BWP7T $T=620360 272600 1 0 $X=620070 $Y=268390
X1235 315 379 133 377 316 5 4 AOI22D0BWP7T $T=621480 335320 1 0 $X=621190 $Y=331110
X1236 320 386 378 382 315 5 4 AOI22D0BWP7T $T=631000 311800 0 180 $X=627350 $Y=307590
X1237 382 387 146 315 316 5 4 AOI22D0BWP7T $T=631560 319640 0 180 $X=627910 $Y=315430
X1238 302 383 315 378 150 5 4 AOI22D0BWP7T $T=629880 280440 1 0 $X=629590 $Y=276230
X1239 302 397 315 395 153 5 4 AOI22D0BWP7T $T=636600 264760 0 0 $X=636310 $Y=264525
X1240 396 400 151 315 316 5 4 AOI22D0BWP7T $T=642760 319640 0 180 $X=639110 $Y=315430
X1241 320 401 395 396 315 5 4 AOI22D0BWP7T $T=641640 288280 1 0 $X=641350 $Y=284070
X1242 162 407 152 129 156 5 4 AOI22D0BWP7T $T=651160 241240 1 180 $X=647510 $Y=241005
X1243 414 409 172 315 156 5 4 AOI22D0BWP7T $T=664040 303960 0 180 $X=660390 $Y=299750
X1244 164 417 315 420 422 5 4 AOI22D0BWP7T $T=665720 303960 1 0 $X=665430 $Y=299750
X1245 180 421 174 129 156 5 4 AOI22D0BWP7T $T=669640 264760 1 180 $X=665990 $Y=264525
X1246 420 426 166 315 156 5 4 AOI22D0BWP7T $T=671320 327480 0 180 $X=667670 $Y=323270
X1247 428 419 182 315 156 5 4 AOI22D0BWP7T $T=673000 280440 0 180 $X=669350 $Y=276230
X1248 168 425 315 183 429 5 4 AOI22D0BWP7T $T=676360 351000 0 180 $X=672710 $Y=346790
X1249 184 430 315 429 433 5 4 AOI22D0BWP7T $T=674680 335320 1 0 $X=674390 $Y=331110
X1250 164 432 315 414 436 5 4 AOI22D0BWP7T $T=676360 280440 1 0 $X=676070 $Y=276230
X1251 184 439 315 406 441 5 4 AOI22D0BWP7T $T=682520 335320 0 0 $X=682230 $Y=335085
X1252 175 440 315 436 453 5 4 AOI22D0BWP7T $T=684200 280440 0 0 $X=683910 $Y=280205
X1253 164 438 315 428 444 5 4 AOI22D0BWP7T $T=685320 272600 0 0 $X=685030 $Y=272365
X1254 168 443 315 189 406 5 4 AOI22D0BWP7T $T=690360 343160 1 180 $X=686710 $Y=342925
X1255 175 447 315 422 452 5 4 AOI22D0BWP7T $T=691480 280440 1 0 $X=691190 $Y=276230
X1256 164 450 129 194 196 5 4 AOI22D0BWP7T $T=693160 241240 0 0 $X=692870 $Y=241005
X1257 175 454 129 444 449 5 4 AOI22D0BWP7T $T=696520 272600 0 180 $X=692870 $Y=268390
X1258 171 451 315 453 456 5 4 AOI22D0BWP7T $T=693160 288280 1 0 $X=692870 $Y=284070
X1259 167 457 315 456 471 5 4 AOI22D0BWP7T $T=702680 296120 0 0 $X=702390 $Y=295885
X1260 168 462 198 199 472 5 4 AOI22D0BWP7T $T=713320 351000 1 0 $X=713030 $Y=346790
X1261 163 476 315 471 477 5 4 AOI22D0BWP7T $T=717240 303960 1 0 $X=716950 $Y=299750
X1262 184 468 198 472 470 5 4 AOI22D0BWP7T $T=720600 343160 0 180 $X=716950 $Y=338950
X1263 168 479 198 202 481 5 4 AOI22D0BWP7T $T=720600 351000 0 0 $X=720310 $Y=350765
X1264 171 464 315 452 475 5 4 AOI22D0BWP7T $T=721720 280440 0 0 $X=721430 $Y=280205
X1265 171 473 129 449 474 5 4 AOI22D0BWP7T $T=722840 256920 1 0 $X=722550 $Y=252710
X1266 184 486 198 481 487 5 4 AOI22D0BWP7T $T=725080 343160 0 0 $X=724790 $Y=342925
X1267 167 485 315 475 488 5 4 AOI22D0BWP7T $T=725640 288280 1 0 $X=725350 $Y=284070
X1268 167 480 129 474 200 5 4 AOI22D0BWP7T $T=735160 249080 0 0 $X=734870 $Y=248845
X1269 163 495 315 488 489 5 4 AOI22D0BWP7T $T=735160 288280 0 0 $X=734870 $Y=288045
X1270 4 5 ICV_41 $T=450120 280440 1 0 $X=449830 $Y=276230
X1271 4 5 ICV_41 $T=477560 343160 1 0 $X=477270 $Y=338950
X1272 4 5 ICV_41 $T=492120 249080 0 0 $X=491830 $Y=248845
X1273 4 5 ICV_41 $T=534120 264760 0 0 $X=533830 $Y=264525
X1274 4 5 ICV_41 $T=534120 311800 1 0 $X=533830 $Y=307590
X1275 4 5 ICV_41 $T=545880 256920 0 0 $X=545590 $Y=256685
X1276 4 5 ICV_41 $T=561560 264760 1 0 $X=561270 $Y=260550
X1277 4 5 ICV_41 $T=576120 296120 1 0 $X=575830 $Y=291910
X1278 4 5 ICV_41 $T=602440 249080 1 0 $X=602150 $Y=244870
X1279 4 5 ICV_41 $T=618120 288280 0 0 $X=617830 $Y=288045
X1280 4 5 ICV_41 $T=618120 351000 1 0 $X=617830 $Y=346790
X1281 4 5 ICV_41 $T=634360 241240 0 0 $X=634070 $Y=241005
X1282 4 5 ICV_41 $T=643880 343160 0 0 $X=643590 $Y=342925
X1283 4 5 ICV_41 $T=644440 358840 1 0 $X=644150 $Y=354630
X1284 4 5 ICV_41 $T=660120 335320 1 0 $X=659830 $Y=331110
X1285 4 5 ICV_41 $T=702120 288280 0 0 $X=701830 $Y=288045
X1286 4 5 ICV_41 $T=720040 264760 0 0 $X=719750 $Y=264525
X1287 4 5 ICV_41 $T=727880 241240 0 0 $X=727590 $Y=241005
X1288 4 5 ICV_41 $T=727880 272600 1 0 $X=727590 $Y=268390
X1289 4 5 ICV_41 $T=729000 319640 0 0 $X=728710 $Y=319405
X1290 4 5 ICV_41 $T=729000 335320 1 0 $X=728710 $Y=331110
X1291 4 5 ICV_37 $T=450120 272600 0 0 $X=449830 $Y=272365
X1292 4 5 ICV_37 $T=470280 343160 1 0 $X=469990 $Y=338950
X1293 4 5 ICV_37 $T=492120 280440 0 0 $X=491830 $Y=280205
X1294 4 5 ICV_37 $T=492120 343160 0 0 $X=491830 $Y=342925
X1295 4 5 ICV_37 $T=501080 319640 0 0 $X=500790 $Y=319405
X1296 4 5 ICV_37 $T=504440 280440 1 0 $X=504150 $Y=276230
X1297 4 5 ICV_37 $T=522920 280440 1 0 $X=522630 $Y=276230
X1298 4 5 ICV_37 $T=529640 343160 1 0 $X=529350 $Y=338950
X1299 4 5 ICV_37 $T=534120 335320 1 0 $X=533830 $Y=331110
X1300 4 5 ICV_37 $T=534120 358840 1 0 $X=533830 $Y=354630
X1301 4 5 ICV_37 $T=547560 249080 1 0 $X=547270 $Y=244870
X1302 4 5 ICV_37 $T=555400 280440 0 0 $X=555110 $Y=280205
X1303 4 5 ICV_37 $T=557080 319640 0 0 $X=556790 $Y=319405
X1304 4 5 ICV_37 $T=571640 249080 0 0 $X=571350 $Y=248845
X1305 4 5 ICV_37 $T=593480 303960 1 0 $X=593190 $Y=299750
X1306 4 5 ICV_37 $T=605240 335320 1 0 $X=604950 $Y=331110
X1307 4 5 ICV_37 $T=618120 335320 1 0 $X=617830 $Y=331110
X1308 4 5 ICV_37 $T=633240 280440 1 0 $X=632950 $Y=276230
X1309 4 5 ICV_37 $T=638840 351000 0 0 $X=638550 $Y=350765
X1310 4 5 ICV_37 $T=647240 272600 1 0 $X=646950 $Y=268390
X1311 4 5 ICV_37 $T=655640 272600 0 0 $X=655350 $Y=272365
X1312 4 5 ICV_37 $T=655640 311800 1 0 $X=655350 $Y=307590
X1313 4 5 ICV_37 $T=655640 327480 0 0 $X=655350 $Y=327245
X1314 4 5 ICV_37 $T=660120 264760 1 0 $X=659830 $Y=260550
X1315 4 5 ICV_37 $T=662920 351000 0 0 $X=662630 $Y=350765
X1316 4 5 ICV_37 $T=673000 280440 1 0 $X=672710 $Y=276230
X1317 4 5 ICV_37 $T=697640 272600 0 0 $X=697350 $Y=272365
X1318 4 5 ICV_37 $T=724520 272600 0 0 $X=724230 $Y=272365
X1319 4 5 ICV_43 $T=450120 272600 1 0 $X=449830 $Y=268390
X1320 4 5 ICV_43 $T=450120 303960 0 0 $X=449830 $Y=303725
X1321 4 5 ICV_43 $T=496040 296120 1 0 $X=495750 $Y=291910
X1322 4 5 ICV_43 $T=496040 319640 1 0 $X=495750 $Y=315430
X1323 4 5 ICV_43 $T=534120 249080 1 0 $X=533830 $Y=244870
X1324 4 5 ICV_43 $T=534120 288280 1 0 $X=533830 $Y=284070
X1325 4 5 ICV_43 $T=534120 288280 0 0 $X=533830 $Y=288045
X1326 4 5 ICV_43 $T=576120 256920 0 0 $X=575830 $Y=256685
X1327 4 5 ICV_43 $T=593480 311800 0 0 $X=593190 $Y=311565
X1328 4 5 ICV_43 $T=597960 249080 0 0 $X=597670 $Y=248845
X1329 4 5 ICV_43 $T=599640 288280 0 0 $X=599350 $Y=288045
X1330 4 5 ICV_43 $T=600200 303960 0 0 $X=599910 $Y=303725
X1331 4 5 ICV_43 $T=627080 280440 1 0 $X=626790 $Y=276230
X1332 4 5 ICV_43 $T=639960 327480 1 0 $X=639670 $Y=323270
X1333 4 5 ICV_43 $T=660120 343160 1 0 $X=659830 $Y=338950
X1334 4 5 ICV_43 $T=682520 272600 0 0 $X=682230 $Y=272365
X1335 4 5 ICV_43 $T=688680 280440 1 0 $X=688390 $Y=276230
X1336 4 5 ICV_43 $T=690360 241240 0 0 $X=690070 $Y=241005
X1337 4 5 ICV_43 $T=702120 272600 0 0 $X=701830 $Y=272365
X1338 4 5 ICV_43 $T=720040 303960 0 0 $X=719750 $Y=303725
X1339 4 5 ICV_52 $T=450120 335320 1 0 $X=449830 $Y=331110
X1340 4 5 ICV_52 $T=459080 296120 1 0 $X=458790 $Y=291910
X1341 4 5 ICV_52 $T=475880 280440 1 0 $X=475590 $Y=276230
X1342 4 5 ICV_52 $T=492120 358840 1 0 $X=491830 $Y=354630
X1343 4 5 ICV_52 $T=501080 241240 0 0 $X=500790 $Y=241005
X1344 4 5 ICV_52 $T=529080 256920 0 0 $X=528790 $Y=256685
X1345 4 5 ICV_52 $T=543080 335320 0 0 $X=542790 $Y=335085
X1346 4 5 ICV_52 $T=547000 319640 0 0 $X=546710 $Y=319405
X1347 4 5 ICV_52 $T=550920 296120 0 0 $X=550630 $Y=295885
X1348 4 5 ICV_52 $T=559880 319640 1 0 $X=559590 $Y=315430
X1349 4 5 ICV_52 $T=561000 296120 1 0 $X=560710 $Y=291910
X1350 4 5 ICV_52 $T=576120 288280 1 0 $X=575830 $Y=284070
X1351 4 5 ICV_52 $T=603000 256920 1 0 $X=602710 $Y=252710
X1352 4 5 ICV_52 $T=605240 272600 0 0 $X=604950 $Y=272365
X1353 4 5 ICV_52 $T=605800 343160 1 0 $X=605510 $Y=338950
X1354 4 5 ICV_52 $T=613080 288280 1 0 $X=612790 $Y=284070
X1355 4 5 ICV_52 $T=648360 264760 1 0 $X=648070 $Y=260550
X1356 4 5 ICV_52 $T=655080 296120 1 0 $X=654790 $Y=291910
X1357 4 5 ICV_52 $T=660120 358840 1 0 $X=659830 $Y=354630
X1358 4 5 ICV_52 $T=669080 351000 1 0 $X=668790 $Y=346790
X1359 4 5 ICV_52 $T=705480 343160 1 0 $X=705190 $Y=338950
X1360 4 5 ICV_52 $T=723960 296120 0 0 $X=723670 $Y=295885
X1361 4 5 ICV_52 $T=723960 311800 0 0 $X=723670 $Y=311565
X1362 4 5 ICV_38 $T=486520 327480 0 0 $X=486230 $Y=327245
X1363 4 5 ICV_38 $T=486520 351000 1 0 $X=486230 $Y=346790
X1364 4 5 ICV_38 $T=528520 249080 1 0 $X=528230 $Y=244870
X1365 4 5 ICV_38 $T=528520 264760 1 0 $X=528230 $Y=260550
X1366 4 5 ICV_38 $T=528520 280440 1 0 $X=528230 $Y=276230
X1367 4 5 ICV_38 $T=528520 319640 0 0 $X=528230 $Y=319405
X1368 4 5 ICV_38 $T=528520 327480 1 0 $X=528230 $Y=323270
X1369 4 5 ICV_38 $T=612520 296120 1 0 $X=612230 $Y=291910
X1370 4 5 ICV_38 $T=612520 303960 1 0 $X=612230 $Y=299750
X1371 4 5 ICV_38 $T=612520 311800 1 0 $X=612230 $Y=307590
X1372 4 5 ICV_38 $T=654520 241240 0 0 $X=654230 $Y=241005
X1373 4 5 ICV_38 $T=654520 264760 1 0 $X=654230 $Y=260550
X1374 4 5 ICV_38 $T=654520 272600 1 0 $X=654230 $Y=268390
X1375 4 5 ICV_38 $T=654520 311800 0 0 $X=654230 $Y=311565
X1376 4 5 ICV_38 $T=696520 256920 0 0 $X=696230 $Y=256685
X1377 4 5 ICV_38 $T=696520 272600 1 0 $X=696230 $Y=268390
X1378 4 5 ICV_38 $T=696520 280440 0 0 $X=696230 $Y=280205
X1379 4 5 ICV_38 $T=696520 288280 1 0 $X=696230 $Y=284070
X1380 4 5 ICV_38 $T=696520 327480 1 0 $X=696230 $Y=323270
X1381 4 5 ICV_38 $T=696520 335320 0 0 $X=696230 $Y=335085
X1382 4 5 ICV_38 $T=696520 358840 1 0 $X=696230 $Y=354630
X1383 4 5 ICV_45 $T=461320 351000 0 0 $X=461030 $Y=350765
X1384 4 5 ICV_45 $T=462440 327480 1 0 $X=462150 $Y=323270
X1385 4 5 ICV_45 $T=463000 256920 0 0 $X=462710 $Y=256685
X1386 4 5 ICV_45 $T=502200 256920 0 0 $X=501910 $Y=256685
X1387 4 5 ICV_45 $T=506120 280440 0 0 $X=505830 $Y=280205
X1388 4 5 ICV_45 $T=534120 296120 1 0 $X=533830 $Y=291910
X1389 4 5 ICV_45 $T=545880 311800 0 0 $X=545590 $Y=311565
X1390 4 5 ICV_45 $T=546440 327480 1 0 $X=546150 $Y=323270
X1391 4 5 ICV_45 $T=547000 343160 1 0 $X=546710 $Y=338950
X1392 4 5 ICV_45 $T=576120 256920 1 0 $X=575830 $Y=252710
X1393 4 5 ICV_45 $T=581720 311800 1 0 $X=581430 $Y=307590
X1394 4 5 ICV_45 $T=589560 351000 1 0 $X=589270 $Y=346790
X1395 4 5 ICV_45 $T=660120 249080 1 0 $X=659830 $Y=244870
X1396 4 5 ICV_45 $T=660120 256920 0 0 $X=659830 $Y=256685
X1397 4 5 ICV_45 $T=660120 272600 1 0 $X=659830 $Y=268390
X1398 4 5 ICV_45 $T=660120 296120 1 0 $X=659830 $Y=291910
X1399 4 5 ICV_45 $T=660120 296120 0 0 $X=659830 $Y=295885
X1400 4 5 ICV_45 $T=672440 327480 0 0 $X=672150 $Y=327245
X1401 4 5 ICV_45 $T=713880 335320 0 0 $X=713590 $Y=335085
X1402 391 4 5 398 BUFFD3BWP7T $T=635480 351000 1 0 $X=635190 $Y=346790
X1403 177 4 5 74 BUFFD3BWP7T $T=666280 249080 1 180 $X=662070 $Y=248845
X1404 366 4 5 391 BUFFD1BWP7T $T=631560 351000 1 0 $X=631270 $Y=346790
X1405 374 4 5 408 BUFFD1BWP7T $T=660680 343160 0 0 $X=660390 $Y=342925
X1406 27 16 4 5 INVD12BWP7T $T=460200 319640 0 180 $X=450390 $Y=315430
X1407 16 5 7 4 CKND12BWP7T $T=463000 335320 0 180 $X=453750 $Y=331110
X1408 16 5 58 4 CKND12BWP7T $T=543640 264760 0 180 $X=534390 $Y=260550
X1409 16 5 149 4 CKND12BWP7T $T=687560 256920 0 0 $X=687270 $Y=256685
X1410 58 301 104 4 5 DFQD2BWP7T $T=553160 311800 1 0 $X=552870 $Y=307590
X1411 149 413 182 4 5 DFQD2BWP7T $T=661240 288280 0 0 $X=660950 $Y=288045
X1412 149 412 172 4 5 DFQD2BWP7T $T=673000 311800 1 180 $X=661510 $Y=311565
X1413 19 4 5 129 BUFFD5BWP7T $T=591800 249080 0 0 $X=591510 $Y=248845
X1414 19 4 5 315 BUFFD5BWP7T $T=608600 288280 1 180 $X=602150 $Y=288045
X1415 140 145 4 5 BUFFD2BWP7T $T=622600 343160 0 0 $X=622310 $Y=342925
X1416 191 85 4 5 BUFFD2BWP7T $T=690920 296120 1 180 $X=687270 $Y=295885
X1417 79 80 296 4 5 ND2D2BWP7T $T=540280 327480 1 180 $X=536070 $Y=327245
X1418 92 336 341 4 5 ND2D2BWP7T $T=585640 335320 1 0 $X=585350 $Y=331110
X1419 336 106 385 4 5 ND2D2BWP7T $T=629320 272600 1 0 $X=629030 $Y=268390
X1420 336 118 45 4 5 ND2D2BWP7T $T=647240 272600 0 180 $X=643030 $Y=268390
X1421 336 116 79 4 5 ND2D2BWP7T $T=643880 256920 0 0 $X=643590 $Y=256685
X1422 79 163 398 4 5 ND2D2BWP7T $T=648360 288280 1 0 $X=648070 $Y=284070
X1423 408 167 398 4 5 ND2D2BWP7T $T=649480 296120 0 0 $X=649190 $Y=295885
X1424 45 171 398 4 5 ND2D2BWP7T $T=650600 272600 1 0 $X=650310 $Y=268390
X1425 83 4 79 11 5 CKND2D2BWP7T $T=541400 358840 0 180 $X=537190 $Y=354630
X1426 76 4 82 98 5 CKND2D2BWP7T $T=558200 241240 1 180 $X=553990 $Y=241005
X1427 45 10 43 4 5 ND2D1P5BWP7T $T=476440 303960 1 0 $X=476150 $Y=299750
X1428 60 37 43 4 5 ND2D1P5BWP7T $T=506120 303960 1 180 $X=501910 $Y=303725
X1429 79 50 43 4 5 ND2D1P5BWP7T $T=538600 311800 1 180 $X=534390 $Y=311565
X1430 77 81 76 4 5 ND2D1P5BWP7T $T=540840 249080 0 180 $X=536630 $Y=244870
X1431 91 59 93 4 5 ND2D1P5BWP7T $T=550920 358840 0 180 $X=546710 $Y=354630
X1432 69 94 76 4 5 ND2D1P5BWP7T $T=549240 311800 1 0 $X=548950 $Y=307590
X1433 300 97 95 4 5 ND2D1P5BWP7T $T=556520 256920 0 180 $X=552310 $Y=252710
X1434 336 302 120 4 5 ND2D1P5BWP7T $T=583960 288280 0 180 $X=579750 $Y=284070
X1435 336 316 147 4 5 ND2D1P5BWP7T $T=625960 351000 0 0 $X=625670 $Y=350765
X1436 155 320 336 4 5 ND2D1P5BWP7T $T=646120 351000 1 180 $X=641910 $Y=350765
X1437 145 156 398 4 5 ND2D1P5BWP7T $T=642760 327480 1 0 $X=642470 $Y=323270
X1438 159 164 398 4 5 ND2D1P5BWP7T $T=648360 311800 0 0 $X=648070 $Y=311565
X1439 385 168 161 4 5 ND2D1P5BWP7T $T=650040 351000 0 0 $X=649750 $Y=350765
X1440 144 175 398 4 5 ND2D1P5BWP7T $T=660680 280440 1 0 $X=660390 $Y=276230
X1441 4 5 ICV_64 $T=485960 280440 0 0 $X=485670 $Y=280205
X1442 4 5 ICV_64 $T=485960 303960 0 0 $X=485670 $Y=303725
X1443 4 5 ICV_64 $T=485960 311800 0 0 $X=485670 $Y=311565
X1444 4 5 ICV_64 $T=527960 249080 0 0 $X=527670 $Y=248845
X1445 4 5 ICV_64 $T=527960 288280 0 0 $X=527670 $Y=288045
X1446 4 5 ICV_64 $T=527960 311800 1 0 $X=527670 $Y=307590
X1447 4 5 ICV_64 $T=527960 335320 0 0 $X=527670 $Y=335085
X1448 4 5 ICV_64 $T=527960 351000 1 0 $X=527670 $Y=346790
X1449 4 5 ICV_64 $T=569960 319640 0 0 $X=569670 $Y=319405
X1450 4 5 ICV_64 $T=569960 335320 1 0 $X=569670 $Y=331110
X1451 4 5 ICV_64 $T=569960 343160 0 0 $X=569670 $Y=342925
X1452 4 5 ICV_64 $T=569960 351000 0 0 $X=569670 $Y=350765
X1453 4 5 ICV_64 $T=611960 256920 0 0 $X=611670 $Y=256685
X1454 4 5 ICV_64 $T=611960 343160 1 0 $X=611670 $Y=338950
X1455 4 5 ICV_64 $T=611960 351000 0 0 $X=611670 $Y=350765
X1456 4 5 ICV_64 $T=653960 280440 0 0 $X=653670 $Y=280205
X1457 4 5 ICV_64 $T=653960 303960 0 0 $X=653670 $Y=303725
X1458 4 5 ICV_64 $T=653960 335320 0 0 $X=653670 $Y=335085
X1459 4 5 ICV_64 $T=653960 343160 1 0 $X=653670 $Y=338950
X1460 4 5 ICV_64 $T=653960 351000 0 0 $X=653670 $Y=350765
X1461 4 5 ICV_64 $T=695960 264760 0 0 $X=695670 $Y=264525
X1462 4 5 ICV_64 $T=695960 303960 0 0 $X=695670 $Y=303725
X1463 4 5 ICV_64 $T=695960 319640 0 0 $X=695670 $Y=319405
X1464 4 5 ICV_64 $T=737960 280440 1 0 $X=737670 $Y=276230
X1465 4 5 ICV_64 $T=737960 288280 1 0 $X=737670 $Y=284070
X1466 4 5 ICV_64 $T=737960 327480 0 0 $X=737670 $Y=327245
X1467 124 123 5 122 121 4 IAO21D1BWP7T $T=589560 351000 0 180 $X=585350 $Y=346790
X1468 90 89 5 92 296 4 OAI21D1BWP7T $T=548680 327480 0 0 $X=548390 $Y=327245
X1469 184 188 5 439 399 4 OAI21D1BWP7T $T=681400 343160 0 0 $X=681110 $Y=342925
X1528 43 291 267 4 5 INR2XD2BWP7T $T=539720 311800 0 0 $X=539430 $Y=311565
X1529 336 126 125 4 5 INR2XD2BWP7T $T=595160 288280 0 180 $X=588710 $Y=284070
X1530 398 158 169 4 5 INR2XD2BWP7T $T=653960 343160 0 180 $X=647510 $Y=338950
X1531 4 5 ICV_66 $T=450120 288280 0 0 $X=449830 $Y=288045
X1532 4 5 ICV_66 $T=468040 311800 1 0 $X=467750 $Y=307590
X1533 4 5 ICV_66 $T=468040 319640 0 0 $X=467750 $Y=319405
X1534 4 5 ICV_66 $T=502200 351000 0 0 $X=501910 $Y=350765
X1535 4 5 ICV_66 $T=503320 249080 1 0 $X=503030 $Y=244870
X1536 4 5 ICV_66 $T=509480 272600 1 0 $X=509190 $Y=268390
X1537 4 5 ICV_66 $T=509480 296120 1 0 $X=509190 $Y=291910
X1538 4 5 ICV_66 $T=509480 319640 1 0 $X=509190 $Y=315430
X1539 4 5 ICV_66 $T=552040 327480 0 0 $X=551750 $Y=327245
X1540 4 5 ICV_66 $T=552040 335320 0 0 $X=551750 $Y=335085
X1541 4 5 ICV_66 $T=576120 327480 0 0 $X=575830 $Y=327245
X1542 4 5 ICV_66 $T=594040 296120 0 0 $X=593750 $Y=295885
X1543 4 5 ICV_66 $T=594040 335320 0 0 $X=593750 $Y=335085
X1544 4 5 ICV_66 $T=618120 296120 1 0 $X=617830 $Y=291910
X1545 4 5 ICV_66 $T=634920 256920 1 0 $X=634630 $Y=252710
X1546 4 5 ICV_66 $T=660120 256920 1 0 $X=659830 $Y=252710
X1547 4 5 ICV_66 $T=660120 280440 0 0 $X=659830 $Y=280205
X1548 4 5 ICV_66 $T=678040 335320 1 0 $X=677750 $Y=331110
X1549 4 5 ICV_66 $T=702120 249080 1 0 $X=701830 $Y=244870
X1550 4 5 7 214 8 ICV_65 $T=450120 327480 1 0 $X=449830 $Y=323270
X1551 4 5 7 223 28 ICV_65 $T=459080 351000 1 0 $X=458790 $Y=346790
X1552 4 5 7 227 217 ICV_65 $T=463000 335320 1 0 $X=462710 $Y=331110
X1553 4 5 13 226 221 ICV_65 $T=463560 280440 1 0 $X=463270 $Y=276230
X1554 4 5 7 232 228 ICV_65 $T=470840 343160 0 0 $X=470550 $Y=342925
X1555 4 5 13 237 3 ICV_65 $T=472520 288280 0 0 $X=472230 $Y=288045
X1556 4 5 7 239 231 ICV_65 $T=473640 303960 0 0 $X=473350 $Y=303725
X1557 4 5 58 271 251 ICV_65 $T=508360 264760 1 0 $X=508070 $Y=260550
X1558 4 5 58 280 244 ICV_65 $T=510040 272600 0 0 $X=509750 $Y=272365
X1559 4 5 58 283 264 ICV_65 $T=511720 288280 0 0 $X=511430 $Y=288045
X1560 4 5 58 294 247 ICV_65 $T=534120 272600 0 0 $X=533830 $Y=272365
X1561 4 5 58 337 333 ICV_65 $T=581720 296120 0 0 $X=581430 $Y=295885
X1562 4 5 149 389 382 ICV_65 $T=622600 303960 1 0 $X=622310 $Y=299750
X1563 4 5 149 404 396 ICV_65 $T=634920 303960 1 0 $X=634630 $Y=299750
X1564 4 5 149 437 420 ICV_65 $T=673000 311800 0 0 $X=672710 $Y=311565
X1565 4 5 149 467 444 ICV_65 $T=702120 264760 1 0 $X=701830 $Y=260550
X1566 4 5 149 455 453 ICV_65 $T=702120 288280 1 0 $X=701830 $Y=284070
X1567 4 5 149 482 475 ICV_65 $T=715560 288280 0 0 $X=715270 $Y=288045
X1568 19 24 4 5 BUFFD4BWP7T $T=455160 288280 1 0 $X=454870 $Y=284070
X1569 4 5 ICV_51 $T=489320 241240 0 0 $X=489030 $Y=241005
X1570 4 5 ICV_51 $T=489320 288280 0 0 $X=489030 $Y=288045
X1571 4 5 ICV_51 $T=489320 296120 1 0 $X=489030 $Y=291910
X1572 4 5 ICV_51 $T=489320 303960 1 0 $X=489030 $Y=299750
X1573 4 5 ICV_51 $T=489320 327480 1 0 $X=489030 $Y=323270
X1574 4 5 ICV_51 $T=531320 241240 0 0 $X=531030 $Y=241005
X1575 4 5 ICV_51 $T=531320 272600 0 0 $X=531030 $Y=272365
X1576 4 5 ICV_51 $T=531320 311800 0 0 $X=531030 $Y=311565
X1577 4 5 ICV_51 $T=531320 343160 0 0 $X=531030 $Y=342925
X1578 4 5 ICV_51 $T=573320 256920 1 0 $X=573030 $Y=252710
X1579 4 5 ICV_51 $T=573320 311800 1 0 $X=573030 $Y=307590
X1580 4 5 ICV_51 $T=573320 327480 1 0 $X=573030 $Y=323270
X1581 4 5 ICV_51 $T=615320 280440 0 0 $X=615030 $Y=280205
X1582 4 5 ICV_51 $T=615320 288280 0 0 $X=615030 $Y=288045
X1583 4 5 ICV_51 $T=615320 335320 1 0 $X=615030 $Y=331110
X1584 4 5 ICV_51 $T=615320 343160 0 0 $X=615030 $Y=342925
X1585 4 5 ICV_51 $T=657320 249080 1 0 $X=657030 $Y=244870
X1586 4 5 ICV_51 $T=657320 256920 1 0 $X=657030 $Y=252710
X1587 4 5 ICV_51 $T=657320 319640 0 0 $X=657030 $Y=319405
X1588 4 5 ICV_51 $T=657320 343160 0 0 $X=657030 $Y=342925
X1589 4 5 ICV_51 $T=657320 351000 1 0 $X=657030 $Y=346790
X1590 4 5 ICV_51 $T=699320 249080 0 0 $X=699030 $Y=248845
X1591 4 5 ICV_51 $T=699320 264760 1 0 $X=699030 $Y=260550
X1592 4 5 ICV_51 $T=699320 288280 0 0 $X=699030 $Y=288045
X1593 4 5 ICV_51 $T=699320 303960 1 0 $X=699030 $Y=299750
X1594 4 5 ICV_51 $T=699320 319640 1 0 $X=699030 $Y=315430
X1595 4 5 ICV_51 $T=699320 327480 0 0 $X=699030 $Y=327245
X1596 4 5 ICV_51 $T=699320 343160 0 0 $X=699030 $Y=342925
X1597 4 5 ICV_51 $T=699320 351000 0 0 $X=699030 $Y=350765
X1598 92 4 88 90 89 5 OAI21D2BWP7T $T=552040 335320 1 180 $X=546710 $Y=335085
X1599 89 5 90 102 4 76 NR3D3BWP7T $T=552600 343160 0 0 $X=552310 $Y=342925
X1600 89 103 102 101 5 4 292 OR4D1BWP7T $T=564920 358840 0 180 $X=560150 $Y=354630
X1601 89 102 109 107 5 4 305 OR4D1BWP7T $T=569960 343160 1 180 $X=565190 $Y=342925
X1602 89 4 109 103 5 335 IND3D0BWP7T $T=576680 351000 1 0 $X=576390 $Y=346790
X1603 89 4 109 103 5 341 IND3D0BWP7T $T=582280 351000 1 0 $X=581990 $Y=346790
X1604 124 123 122 291 5 4 IAO21D2BWP7T $T=600760 343160 1 180 $X=595430 $Y=342925
X1605 137 124 139 92 4 5 393 OA31D0BWP7T $T=629880 358840 1 0 $X=629590 $Y=354630
.ENDS
***************************************
.SUBCKT ICV_59
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_62
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_39 1 2
** N=2 EP=2 IP=4 FDC=6
*.SEEDPROM
X1 1 2 ICV_38 $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_42 1 2
** N=2 EP=2 IP=4 FDC=22
*.SEEDPROM
X0 1 2 ICV_40 $T=8960 0 0 0 $X=8670 $Y=-235
X1 1 2 DCAP16BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT OA32D0BWP7T A1 A2 A3 B2 B1 VDD VSS Z
** N=13 EP=8 IP=0 FDC=12
*.SEEDPROM
M0 9 A1 10 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=750 $D=0
M1 10 A2 9 VSS N L=1.8e-07 W=5e-07 $X=1340 $Y=750 $D=0
M2 9 A3 10 VSS N L=1.8e-07 W=5e-07 $X=2060 $Y=750 $D=0
M3 VSS B2 9 VSS N L=1.8e-07 W=5e-07 $X=2780 $Y=750 $D=0
M4 9 B1 VSS VSS N L=1.8e-07 W=5e-07 $X=3500 $Y=750 $D=0
M5 Z 10 VSS VSS N L=1.8e-07 W=4.65e-07 $X=4760 $Y=880 $D=0
M6 11 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2860 $D=16
M7 12 A2 11 VDD P L=1.8e-07 W=6.85e-07 $X=1270 $Y=2860 $D=16
M8 10 A3 12 VDD P L=1.8e-07 W=6.85e-07 $X=1920 $Y=2860 $D=16
M9 13 B2 10 VDD P L=1.8e-07 W=6.85e-07 $X=2780 $Y=2860 $D=16
M10 VDD B1 13 VDD P L=1.8e-07 W=6.85e-07 $X=3500 $Y=2860 $D=16
M11 Z 10 VDD VDD P L=1.8e-07 W=6.85e-07 $X=4380 $Y=2860 $D=16
.ENDS
***************************************
.SUBCKT BUFFD6BWP7T I Z VSS VDD
** N=5 EP=4 IP=0 FDC=16
*.SEEDPROM
M0 5 I VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=2080 $Y=345 $D=0
M3 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=2800 $Y=345 $D=0
M4 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=3520 $Y=345 $D=0
M5 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=4240 $Y=345 $D=0
M6 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=4960 $Y=345 $D=0
M7 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=5680 $Y=345 $D=0
M8 5 I VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M9 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M10 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2080 $Y=2205 $D=16
M11 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=2800 $Y=2205 $D=16
M12 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3520 $Y=2205 $D=16
M13 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=4240 $Y=2205 $D=16
M14 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4960 $Y=2205 $D=16
M15 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=5680 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OAI31D2BWP7T B VSS ZN A3 A1 A2 VDD
** N=12 EP=7 IP=0 FDC=16
*.SEEDPROM
M0 VSS B 8 VSS N L=1.8e-07 W=9.3e-07 $X=620 $Y=345 $D=0
M1 8 B VSS VSS N L=1.8e-07 W=9.3e-07 $X=1420 $Y=345 $D=0
M2 ZN A1 8 VSS N L=1.8e-07 W=9.3e-07 $X=2140 $Y=345 $D=0
M3 8 A1 ZN VSS N L=1.8e-07 W=9.3e-07 $X=2860 $Y=345 $D=0
M4 ZN A3 8 VSS N L=1.8e-07 W=9.3e-07 $X=3580 $Y=345 $D=0
M5 8 A3 ZN VSS N L=1.8e-07 W=9.3e-07 $X=4300 $Y=345 $D=0
M6 ZN A2 8 VSS N L=1.8e-07 W=9.3e-07 $X=5020 $Y=345 $D=0
M7 8 A2 ZN VSS N L=1.8e-07 W=9.3e-07 $X=5740 $Y=345 $D=0
M8 ZN B VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M9 VDD B ZN VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M10 9 A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2140 $Y=2205 $D=16
M11 10 A2 9 VDD P L=1.8e-07 W=1.25e-06 $X=2860 $Y=2325 $D=16
M12 ZN A3 10 VDD P L=1.8e-07 W=1.305e-06 $X=3580 $Y=2270 $D=16
M13 11 A3 ZN VDD P L=1.8e-07 W=1.305e-06 $X=4300 $Y=2270 $D=16
M14 12 A2 11 VDD P L=1.8e-07 W=1.25e-06 $X=5020 $Y=2325 $D=16
M15 VDD A1 12 VDD P L=1.8e-07 W=1.25e-06 $X=5740 $Y=2325 $D=16
.ENDS
***************************************
.SUBCKT ND2D3BWP7T A2 VSS ZN A1 VDD
** N=6 EP=5 IP=0 FDC=12
*.SEEDPROM
M0 6 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS A2 6 VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 6 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=2060 $Y=345 $D=0
M3 ZN A1 6 VSS N L=1.8e-07 W=1e-06 $X=2780 $Y=345 $D=0
M4 6 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=3500 $Y=345 $D=0
M5 ZN A1 6 VSS N L=1.8e-07 W=1e-06 $X=4220 $Y=345 $D=0
M6 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M7 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M8 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M9 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M10 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3500 $Y=2205 $D=16
M11 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4220 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKND0BWP7T I VSS VDD ZN
** N=4 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 ZN I VSS VSS N L=1.8e-07 W=4.2e-07 $X=830 $Y=505 $D=0
M1 ZN I VDD VDD P L=1.8e-07 W=1.13e-06 $X=830 $Y=2445 $D=16
.ENDS
***************************************
.SUBCKT AO211D0BWP7T A1 A2 B C VSS VDD Z
** N=11 EP=7 IP=0 FDC=10
*.SEEDPROM
M0 9 A1 8 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=845 $D=0
M1 VSS A2 9 VSS N L=1.8e-07 W=5e-07 $X=1050 $Y=845 $D=0
M2 8 B VSS VSS N L=1.8e-07 W=5e-07 $X=1780 $Y=880 $D=0
M3 VSS C 8 VSS N L=1.8e-07 W=5e-07 $X=2500 $Y=880 $D=0
M4 Z 8 VSS VSS N L=1.8e-07 W=5e-07 $X=3120 $Y=580 $D=0
M5 8 A1 10 VDD P L=1.8e-07 W=6.85e-07 $X=570 $Y=2395 $D=16
M6 10 A2 8 VDD P L=1.8e-07 W=6.85e-07 $X=1290 $Y=2395 $D=16
M7 11 B 10 VDD P L=1.8e-07 W=6.85e-07 $X=1970 $Y=2790 $D=16
M8 VDD C 11 VDD P L=1.8e-07 W=6.85e-07 $X=2400 $Y=2790 $D=16
M9 Z 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=3120 $Y=2790 $D=16
.ENDS
***************************************
.SUBCKT ICV_63 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230
** N=616 EP=229 IP=4748 FDC=11529
*.SEEDPROM
M0 50 27 3 3 N L=1.8e-07 W=5e-07 $X=460820 $Y=482960 $D=0
M1 3 254 50 3 N L=1.8e-07 W=5e-07 $X=461540 $Y=482960 $D=0
M2 254 256 3 3 N L=1.8e-07 W=5e-07 $X=462200 $Y=483280 $D=0
M3 305 94 3 3 N L=1.8e-07 W=1e-06 $X=514770 $Y=435895 $D=0
M4 3 312 65 3 N L=1.8e-07 W=5.7e-07 $X=514870 $Y=445425 $D=0
M5 65 312 3 3 N L=1.8e-07 W=5.7e-07 $X=515590 $Y=445425 $D=0
M6 592 96 305 3 N L=1.8e-07 W=1e-06 $X=515610 $Y=435895 $D=0
M7 3 312 65 3 N L=1.8e-07 W=5.7e-07 $X=516310 $Y=445425 $D=0
M8 593 312 592 3 N L=1.8e-07 W=1e-06 $X=516315 $Y=435895 $D=0
M9 3 303 593 3 N L=1.8e-07 W=1e-06 $X=517020 $Y=435895 $D=0
M10 65 312 3 3 N L=1.8e-07 W=5.7e-07 $X=517030 $Y=445425 $D=0
M11 3 312 65 3 N L=1.8e-07 W=5.7e-07 $X=517750 $Y=445425 $D=0
M12 65 312 3 3 N L=1.8e-07 W=5.7e-07 $X=518470 $Y=445425 $D=0
M13 3 312 65 3 N L=1.8e-07 W=5.7e-07 $X=519190 $Y=445425 $D=0
M14 65 303 3 3 N L=1.8e-07 W=5.7e-07 $X=519910 $Y=445425 $D=0
M15 3 303 65 3 N L=1.8e-07 W=5.7e-07 $X=520630 $Y=445425 $D=0
M16 65 303 3 3 N L=1.8e-07 W=5.7e-07 $X=521350 $Y=445425 $D=0
M17 3 303 65 3 N L=1.8e-07 W=5.7e-07 $X=522070 $Y=445425 $D=0
M18 65 303 3 3 N L=1.8e-07 W=5.7e-07 $X=522790 $Y=445425 $D=0
M19 3 303 65 3 N L=1.8e-07 W=5.7e-07 $X=523510 $Y=445425 $D=0
M20 65 303 3 3 N L=1.8e-07 W=5.7e-07 $X=524230 $Y=445425 $D=0
M21 352 303 3 3 N L=1.8e-07 W=1e-06 $X=538520 $Y=412375 $D=0
M22 3 354 352 3 N L=1.8e-07 W=1e-06 $X=539240 $Y=412375 $D=0
M23 594 358 3 3 N L=1.8e-07 W=5e-07 $X=543160 $Y=453265 $D=0
M24 595 95 594 3 N L=1.8e-07 W=5e-07 $X=543610 $Y=453265 $D=0
M25 362 342 595 3 N L=1.8e-07 W=5e-07 $X=544210 $Y=453640 $D=0
M26 595 345 362 3 N L=1.8e-07 W=5e-07 $X=544930 $Y=453640 $D=0
M27 357 362 3 3 N L=1.8e-07 W=5e-07 $X=546200 $Y=453265 $D=0
M28 374 366 123 3 N L=1.8e-07 W=8e-07 $X=548740 $Y=412470 $D=0
M29 123 366 374 3 N L=1.8e-07 W=8e-07 $X=549460 $Y=412470 $D=0
M30 374 366 123 3 N L=1.8e-07 W=8e-07 $X=550200 $Y=412470 $D=0
M31 3 352 374 3 N L=1.8e-07 W=6e-07 $X=550920 $Y=412670 $D=0
M32 374 352 3 3 N L=1.8e-07 W=6e-07 $X=551640 $Y=412670 $D=0
M33 3 352 374 3 N L=1.8e-07 W=6e-07 $X=552360 $Y=412670 $D=0
M34 3 382 391 3 N L=1.8e-07 W=4.7e-07 $X=560100 $Y=397085 $D=0
M35 391 382 3 3 N L=1.8e-07 W=4.7e-07 $X=560820 $Y=397085 $D=0
M36 3 382 391 3 N L=1.8e-07 W=4.7e-07 $X=561540 $Y=397085 $D=0
M37 391 382 3 3 N L=1.8e-07 W=4.7e-07 $X=562260 $Y=397085 $D=0
M38 596 133 3 3 N L=1.8e-07 W=5e-07 $X=562745 $Y=382705 $D=0
M39 3 382 391 3 N L=1.8e-07 W=4.7e-07 $X=562990 $Y=397085 $D=0
M40 385 392 596 3 N L=1.8e-07 W=5e-07 $X=563355 $Y=383095 $D=0
M41 125 391 3 3 N L=1.8e-07 W=6.1e-07 $X=563710 $Y=397085 $D=0
M42 596 381 385 3 N L=1.8e-07 W=5e-07 $X=564075 $Y=383095 $D=0
M43 3 391 125 3 N L=1.8e-07 W=6.1e-07 $X=564430 $Y=397085 $D=0
M44 3 376 596 3 N L=1.8e-07 W=5e-07 $X=564675 $Y=382840 $D=0
M45 125 391 3 3 N L=1.8e-07 W=6.1e-07 $X=565150 $Y=397085 $D=0
M46 3 391 125 3 N L=1.8e-07 W=6.1e-07 $X=565870 $Y=397085 $D=0
M47 597 354 375 3 N L=1.8e-07 W=1e-06 $X=566100 $Y=421905 $D=0
M48 125 391 3 3 N L=1.8e-07 W=6.1e-07 $X=566600 $Y=397085 $D=0
M49 3 366 597 3 N L=1.8e-07 W=1e-06 $X=566820 $Y=421905 $D=0
M50 3 391 125 3 N L=1.8e-07 W=6.1e-07 $X=567320 $Y=397085 $D=0
M51 125 391 3 3 N L=1.8e-07 W=6.1e-07 $X=568040 $Y=397085 $D=0
M52 598 366 3 3 N L=1.8e-07 W=1e-06 $X=568275 $Y=421905 $D=0
M53 3 391 125 3 N L=1.8e-07 W=6.1e-07 $X=568760 $Y=397085 $D=0
M54 375 401 598 3 N L=1.8e-07 W=1e-06 $X=568995 $Y=421905 $D=0
M55 125 391 3 3 N L=1.8e-07 W=6.1e-07 $X=569480 $Y=397085 $D=0
M56 3 309 375 3 N L=1.8e-07 W=1e-06 $X=569715 $Y=421905 $D=0
M57 3 381 420 3 N L=1.8e-07 W=1e-06 $X=577860 $Y=398385 $D=0
M58 420 381 3 3 N L=1.8e-07 W=1e-06 $X=578660 $Y=398385 $D=0
M59 599 127 420 3 N L=1.8e-07 W=1e-06 $X=579420 $Y=398385 $D=0
M60 3 395 599 3 N L=1.8e-07 W=1e-06 $X=580100 $Y=398385 $D=0
M61 600 395 3 3 N L=1.8e-07 W=1e-06 $X=580900 $Y=398385 $D=0
M62 146 141 3 3 N L=1.8e-07 W=1e-06 $X=581380 $Y=359185 $D=0
M63 420 127 600 3 N L=1.8e-07 W=1e-06 $X=581500 $Y=398385 $D=0
M64 3 94 146 3 N L=1.8e-07 W=1e-06 $X=582100 $Y=359185 $D=0
M65 601 376 3 3 N L=1.8e-07 W=5e-07 $X=582340 $Y=382840 $D=0
M66 146 133 3 3 N L=1.8e-07 W=1e-06 $X=582910 $Y=359185 $D=0
M67 602 130 601 3 N L=1.8e-07 W=5e-07 $X=582930 $Y=382840 $D=0
M68 603 418 420 3 N L=1.8e-07 W=1e-06 $X=583140 $Y=398385 $D=0
M69 392 133 602 3 N L=1.8e-07 W=5e-07 $X=583520 $Y=382840 $D=0
M70 3 130 146 3 N L=1.8e-07 W=1e-06 $X=583630 $Y=359185 $D=0
M71 3 397 603 3 N L=1.8e-07 W=1e-06 $X=583760 $Y=398385 $D=0
M72 3 419 392 3 N L=1.8e-07 W=5e-07 $X=584280 $Y=382840 $D=0
M73 604 397 3 3 N L=1.8e-07 W=1e-06 $X=584560 $Y=398385 $D=0
M74 420 418 604 3 N L=1.8e-07 W=1e-06 $X=585170 $Y=398385 $D=0
M75 94 85 3 3 N L=1.8e-07 W=1e-06 $X=593635 $Y=428055 $D=0
M76 3 85 94 3 N L=1.8e-07 W=1e-06 $X=594355 $Y=428055 $D=0
M77 94 85 3 3 N L=1.8e-07 W=1e-06 $X=595095 $Y=428055 $D=0
M78 3 85 94 3 N L=1.8e-07 W=1e-06 $X=595815 $Y=428055 $D=0
M79 94 85 3 3 N L=1.8e-07 W=1e-06 $X=596555 $Y=428055 $D=0
M80 3 85 94 3 N L=1.8e-07 W=1e-06 $X=597275 $Y=428055 $D=0
M81 94 85 3 3 N L=1.8e-07 W=1e-06 $X=598015 $Y=428055 $D=0
M82 3 85 94 3 N L=1.8e-07 W=1e-06 $X=598735 $Y=428055 $D=0
M83 605 149 433 3 N L=1.8e-07 W=5e-07 $X=619440 $Y=406325 $D=0
M84 3 430 605 3 N L=1.8e-07 W=5e-07 $X=620080 $Y=406325 $D=0
M85 3 141 189 3 N L=1.8e-07 W=6e-07 $X=630710 $Y=429745 $D=0
M86 189 141 3 3 N L=1.8e-07 W=6e-07 $X=631430 $Y=429745 $D=0
M87 3 141 189 3 N L=1.8e-07 W=6e-07 $X=632150 $Y=429745 $D=0
M88 189 141 3 3 N L=1.8e-07 W=6e-07 $X=632870 $Y=429745 $D=0
M89 3 141 189 3 N L=1.8e-07 W=6e-07 $X=633590 $Y=429745 $D=0
M90 189 127 3 3 N L=1.8e-07 W=6e-07 $X=634310 $Y=429745 $D=0
M91 3 127 189 3 N L=1.8e-07 W=6e-07 $X=635030 $Y=429745 $D=0
M92 189 127 3 3 N L=1.8e-07 W=6e-07 $X=635750 $Y=429745 $D=0
M93 3 127 189 3 N L=1.8e-07 W=6e-07 $X=636470 $Y=429745 $D=0
M94 189 127 3 3 N L=1.8e-07 W=6e-07 $X=637190 $Y=429745 $D=0
M95 471 150 469 3 N L=1.8e-07 W=1e-06 $X=637820 $Y=367025 $D=0
M96 3 94 189 3 N L=1.8e-07 W=6e-07 $X=637910 $Y=429745 $D=0
M97 189 94 3 3 N L=1.8e-07 W=6e-07 $X=638630 $Y=429745 $D=0
M98 469 143 471 3 N L=1.8e-07 W=1e-06 $X=638650 $Y=367025 $D=0
M99 3 94 189 3 N L=1.8e-07 W=6e-07 $X=639350 $Y=429745 $D=0
M100 3 124 469 3 N L=1.8e-07 W=1e-06 $X=639560 $Y=367025 $D=0
M101 189 94 3 3 N L=1.8e-07 W=6e-07 $X=640070 $Y=429745 $D=0
M102 180 471 3 3 N L=1.8e-07 W=1e-06 $X=640280 $Y=367025 $D=0
M103 3 94 189 3 N L=1.8e-07 W=6e-07 $X=640790 $Y=429745 $D=0
M104 189 125 3 3 N L=1.8e-07 W=6e-07 $X=641510 $Y=429745 $D=0
M105 3 125 189 3 N L=1.8e-07 W=6e-07 $X=642230 $Y=429745 $D=0
M106 189 125 3 3 N L=1.8e-07 W=6e-07 $X=642950 $Y=429745 $D=0
M107 3 125 189 3 N L=1.8e-07 W=6e-07 $X=643670 $Y=429745 $D=0
M108 189 125 3 3 N L=1.8e-07 W=6e-07 $X=644390 $Y=429745 $D=0
M109 606 27 50 1 P L=1.8e-07 W=1.37e-06 $X=460820 $Y=480705 $D=16
M110 1 254 606 1 P L=1.8e-07 W=1.37e-06 $X=461420 $Y=480705 $D=16
M111 254 256 1 1 P L=1.8e-07 W=6.85e-07 $X=462200 $Y=480705 $D=16
M112 330 94 1 1 P L=1.8e-07 W=1.37e-06 $X=514770 $Y=433665 $D=16
M113 335 312 65 1 P L=1.8e-07 W=1.3e-06 $X=514870 $Y=447355 $D=16
M114 305 96 330 1 P L=1.8e-07 W=1.37e-06 $X=515540 $Y=433665 $D=16
M115 65 312 335 1 P L=1.8e-07 W=1.61e-06 $X=515590 $Y=447045 $D=16
M116 330 312 305 1 P L=1.8e-07 W=1.37e-06 $X=516300 $Y=433665 $D=16
M117 335 312 65 1 P L=1.8e-07 W=1.61e-06 $X=516310 $Y=447045 $D=16
M118 305 303 330 1 P L=1.8e-07 W=1.37e-06 $X=517020 $Y=433665 $D=16
M119 65 312 335 1 P L=1.8e-07 W=1.61e-06 $X=517030 $Y=447045 $D=16
M120 335 312 65 1 P L=1.8e-07 W=1.61e-06 $X=517750 $Y=447045 $D=16
M121 65 312 335 1 P L=1.8e-07 W=1.61e-06 $X=518470 $Y=447045 $D=16
M122 335 312 65 1 P L=1.8e-07 W=1.61e-06 $X=519190 $Y=447045 $D=16
M123 1 303 335 1 P L=1.8e-07 W=1.61e-06 $X=519910 $Y=447045 $D=16
M124 335 303 1 1 P L=1.8e-07 W=1.61e-06 $X=520630 $Y=447045 $D=16
M125 1 303 335 1 P L=1.8e-07 W=1.61e-06 $X=521350 $Y=447045 $D=16
M126 335 303 1 1 P L=1.8e-07 W=1.61e-06 $X=522070 $Y=447045 $D=16
M127 1 303 335 1 P L=1.8e-07 W=1.61e-06 $X=522790 $Y=447045 $D=16
M128 335 303 1 1 P L=1.8e-07 W=1.61e-06 $X=523510 $Y=447045 $D=16
M129 1 303 335 1 P L=1.8e-07 W=1.3e-06 $X=524230 $Y=447355 $D=16
M130 1 303 353 1 P L=1.8e-07 W=1.37e-06 $X=537800 $Y=410145 $D=16
M131 353 303 1 1 P L=1.8e-07 W=1.37e-06 $X=538520 $Y=410145 $D=16
M132 352 354 353 1 P L=1.8e-07 W=1.37e-06 $X=539240 $Y=410145 $D=16
M133 353 354 352 1 P L=1.8e-07 W=1.37e-06 $X=539960 $Y=410145 $D=16
M134 1 358 362 1 P L=1.8e-07 W=6.85e-07 $X=543160 $Y=455810 $D=16
M135 362 95 1 1 P L=1.8e-07 W=6.85e-07 $X=543885 $Y=455810 $D=16
M136 607 342 362 1 P L=1.8e-07 W=6.85e-07 $X=544605 $Y=455810 $D=16
M137 1 345 607 1 P L=1.8e-07 W=6.85e-07 $X=545185 $Y=455810 $D=16
M138 357 362 1 1 P L=1.8e-07 W=6.85e-07 $X=545985 $Y=455810 $D=16
M139 123 366 1 1 P L=1.8e-07 W=1.37e-06 $X=548755 $Y=410145 $D=16
M140 1 366 123 1 P L=1.8e-07 W=1.37e-06 $X=549475 $Y=410145 $D=16
M141 123 366 1 1 P L=1.8e-07 W=1.37e-06 $X=550200 $Y=410145 $D=16
M142 1 352 123 1 P L=1.8e-07 W=1.37e-06 $X=550920 $Y=410145 $D=16
M143 123 352 1 1 P L=1.8e-07 W=1.37e-06 $X=551640 $Y=410145 $D=16
M144 1 352 123 1 P L=1.8e-07 W=1.37e-06 $X=552360 $Y=410145 $D=16
M145 391 382 1 1 P L=1.8e-07 W=1.175e-06 $X=559380 $Y=394465 $D=16
M146 1 382 391 1 P L=1.8e-07 W=1.175e-06 $X=560100 $Y=394465 $D=16
M147 391 382 1 1 P L=1.8e-07 W=1.175e-06 $X=560820 $Y=394465 $D=16
M148 1 382 391 1 P L=1.8e-07 W=1.175e-06 $X=561540 $Y=394465 $D=16
M149 391 382 1 1 P L=1.8e-07 W=1.175e-06 $X=562260 $Y=394465 $D=16
M150 608 392 1 1 P L=1.8e-07 W=6.85e-07 $X=562740 $Y=385250 $D=16
M151 1 382 391 1 P L=1.8e-07 W=1.175e-06 $X=562990 $Y=394465 $D=16
M152 385 381 608 1 P L=1.8e-07 W=6.85e-07 $X=563170 $Y=385250 $D=16
M153 125 391 1 1 P L=1.8e-07 W=1.54e-06 $X=563710 $Y=394465 $D=16
M154 609 133 385 1 P L=1.8e-07 W=6.85e-07 $X=563970 $Y=385250 $D=16
M155 1 391 125 1 P L=1.8e-07 W=1.54e-06 $X=564440 $Y=394465 $D=16
M156 1 376 609 1 P L=1.8e-07 W=6.85e-07 $X=564675 $Y=385250 $D=16
M157 125 391 1 1 P L=1.8e-07 W=1.54e-06 $X=565160 $Y=394465 $D=16
M158 1 391 125 1 P L=1.8e-07 W=1.54e-06 $X=565880 $Y=394465 $D=16
M159 375 354 398 1 P L=1.8e-07 W=1.37e-06 $X=566100 $Y=423765 $D=16
M160 125 391 1 1 P L=1.8e-07 W=1.54e-06 $X=566600 $Y=394465 $D=16
M161 398 366 375 1 P L=1.8e-07 W=1.37e-06 $X=566820 $Y=423765 $D=16
M162 1 391 125 1 P L=1.8e-07 W=1.54e-06 $X=567320 $Y=394465 $D=16
M163 125 391 1 1 P L=1.8e-07 W=1.54e-06 $X=568040 $Y=394465 $D=16
M164 398 366 403 1 P L=1.8e-07 W=1.37e-06 $X=568275 $Y=423765 $D=16
M165 1 391 125 1 P L=1.8e-07 W=1.54e-06 $X=568760 $Y=394465 $D=16
M166 403 401 398 1 P L=1.8e-07 W=1.37e-06 $X=568995 $Y=423765 $D=16
M167 125 391 1 1 P L=1.8e-07 W=1.37e-06 $X=569480 $Y=394465 $D=16
M168 1 309 403 1 P L=1.8e-07 W=1.37e-06 $X=569715 $Y=423765 $D=16
M169 1 381 408 1 P L=1.8e-07 W=1.37e-06 $X=577860 $Y=400245 $D=16
M170 408 381 1 1 P L=1.8e-07 W=1.37e-06 $X=578660 $Y=400245 $D=16
M171 411 127 408 1 P L=1.8e-07 W=1.37e-06 $X=579380 $Y=400245 $D=16
M172 408 395 411 1 P L=1.8e-07 W=1.37e-06 $X=580100 $Y=400245 $D=16
M173 610 94 414 1 P L=1.8e-07 W=1.37e-06 $X=580660 $Y=361045 $D=16
M174 411 395 408 1 P L=1.8e-07 W=1.37e-06 $X=580820 $Y=400245 $D=16
M175 1 141 610 1 P L=1.8e-07 W=1.37e-06 $X=581090 $Y=361045 $D=16
M176 408 127 411 1 P L=1.8e-07 W=1.37e-06 $X=581540 $Y=400245 $D=16
M177 611 141 1 1 P L=1.8e-07 W=1.37e-06 $X=581810 $Y=361045 $D=16
M178 614 376 392 1 P L=1.8e-07 W=6.85e-07 $X=582340 $Y=384610 $D=16
M179 612 94 611 1 P L=1.8e-07 W=1.37e-06 $X=582400 $Y=361045 $D=16
M180 392 130 614 1 P L=1.8e-07 W=6.85e-07 $X=582940 $Y=384610 $D=16
M181 613 133 612 1 P L=1.8e-07 W=1.37e-06 $X=582990 $Y=361045 $D=16
M182 411 418 420 1 P L=1.8e-07 W=1.37e-06 $X=583040 $Y=400245 $D=16
M183 146 130 613 1 P L=1.8e-07 W=1.37e-06 $X=583580 $Y=361045 $D=16
M184 614 133 392 1 P L=1.8e-07 W=6.85e-07 $X=583665 $Y=384610 $D=16
M185 420 397 411 1 P L=1.8e-07 W=1.37e-06 $X=583760 $Y=400245 $D=16
M186 1 419 614 1 P L=1.8e-07 W=6.85e-07 $X=584280 $Y=384610 $D=16
M187 615 130 146 1 P L=1.8e-07 W=1.37e-06 $X=584300 $Y=361045 $D=16
M188 411 397 420 1 P L=1.8e-07 W=1.37e-06 $X=584520 $Y=400245 $D=16
M189 414 133 615 1 P L=1.8e-07 W=1.37e-06 $X=584840 $Y=361045 $D=16
M190 420 418 411 1 P L=1.8e-07 W=1.37e-06 $X=585280 $Y=400245 $D=16
M191 94 85 1 1 P L=1.8e-07 W=1.37e-06 $X=593635 $Y=425825 $D=16
M192 1 85 94 1 P L=1.8e-07 W=1.37e-06 $X=594355 $Y=425825 $D=16
M193 94 85 1 1 P L=1.8e-07 W=1.37e-06 $X=595095 $Y=425825 $D=16
M194 1 85 94 1 P L=1.8e-07 W=1.37e-06 $X=595815 $Y=425825 $D=16
M195 94 85 1 1 P L=1.8e-07 W=1.37e-06 $X=596555 $Y=425825 $D=16
M196 1 85 94 1 P L=1.8e-07 W=1.37e-06 $X=597275 $Y=425825 $D=16
M197 94 85 1 1 P L=1.8e-07 W=1.37e-06 $X=598015 $Y=425825 $D=16
M198 1 85 94 1 P L=1.8e-07 W=1.37e-06 $X=598735 $Y=425825 $D=16
M199 433 149 1 1 P L=1.8e-07 W=6.85e-07 $X=619360 $Y=408510 $D=16
M200 1 430 433 1 P L=1.8e-07 W=6.85e-07 $X=620080 $Y=408510 $D=16
M201 463 141 1 1 P L=1.8e-07 W=1.34e-06 $X=630710 $Y=431635 $D=16
M202 1 141 463 1 P L=1.8e-07 W=1.72e-06 $X=631430 $Y=431255 $D=16
M203 463 141 1 1 P L=1.8e-07 W=1.72e-06 $X=632150 $Y=431255 $D=16
M204 1 141 463 1 P L=1.8e-07 W=1.72e-06 $X=632870 $Y=431255 $D=16
M205 463 141 1 1 P L=1.8e-07 W=1.72e-06 $X=633590 $Y=431255 $D=16
M206 472 127 463 1 P L=1.8e-07 W=1.645e-06 $X=634310 $Y=431330 $D=16
M207 463 127 472 1 P L=1.8e-07 W=1.645e-06 $X=635030 $Y=431330 $D=16
M208 472 127 463 1 P L=1.8e-07 W=1.645e-06 $X=635750 $Y=431330 $D=16
M209 463 127 472 1 P L=1.8e-07 W=1.645e-06 $X=636470 $Y=431330 $D=16
M210 472 127 463 1 P L=1.8e-07 W=1.645e-06 $X=637190 $Y=431330 $D=16
M211 616 150 1 1 P L=1.8e-07 W=1.37e-06 $X=637820 $Y=368885 $D=16
M212 468 94 472 1 P L=1.8e-07 W=1.645e-06 $X=637910 $Y=431330 $D=16
M213 472 94 468 1 P L=1.8e-07 W=1.645e-06 $X=638630 $Y=431330 $D=16
M214 471 143 616 1 P L=1.8e-07 W=1.37e-06 $X=638650 $Y=368885 $D=16
M215 468 94 472 1 P L=1.8e-07 W=1.645e-06 $X=639350 $Y=431330 $D=16
M216 1 124 471 1 P L=1.8e-07 W=1.37e-06 $X=639560 $Y=368885 $D=16
M217 472 94 468 1 P L=1.8e-07 W=1.645e-06 $X=640070 $Y=431330 $D=16
M218 180 471 1 1 P L=1.8e-07 W=1.37e-06 $X=640280 $Y=368885 $D=16
M219 468 94 472 1 P L=1.8e-07 W=1.645e-06 $X=640790 $Y=431330 $D=16
M220 189 125 468 1 P L=1.8e-07 W=1.72e-06 $X=641510 $Y=431255 $D=16
M221 468 125 189 1 P L=1.8e-07 W=1.72e-06 $X=642230 $Y=431255 $D=16
M222 189 125 468 1 P L=1.8e-07 W=1.72e-06 $X=642950 $Y=431255 $D=16
M223 468 125 189 1 P L=1.8e-07 W=1.72e-06 $X=643670 $Y=431255 $D=16
M224 189 125 468 1 P L=1.8e-07 W=1.34e-06 $X=644390 $Y=431635 $D=16
D225 3 382 DN AREA=2.037e-13 PJ=1.81e-06 $X=558900 $Y=396900 $D=32
X244 4 3 PVSS3CDG $T=900240 370000 0 90 $X=780240 $Y=369400
X403 1 3 DCAPBWP7T $T=459080 405880 1 0 $X=458790 $Y=401670
X404 1 3 DCAPBWP7T $T=466920 437240 1 0 $X=466630 $Y=433030
X405 1 3 DCAPBWP7T $T=468600 390200 1 0 $X=468310 $Y=385990
X406 1 3 DCAPBWP7T $T=474200 398040 1 0 $X=473910 $Y=393830
X407 1 3 DCAPBWP7T $T=475880 429400 1 0 $X=475590 $Y=425190
X408 1 3 DCAPBWP7T $T=492120 405880 1 0 $X=491830 $Y=401670
X409 1 3 DCAPBWP7T $T=492120 476440 1 0 $X=491830 $Y=472230
X410 1 3 DCAPBWP7T $T=496600 405880 0 0 $X=496310 $Y=405645
X411 1 3 DCAPBWP7T $T=498840 452920 1 0 $X=498550 $Y=448710
X412 1 3 DCAPBWP7T $T=508920 374520 1 0 $X=508630 $Y=370310
X413 1 3 DCAPBWP7T $T=510040 413720 1 0 $X=509750 $Y=409510
X414 1 3 DCAPBWP7T $T=510040 421560 1 0 $X=509750 $Y=417350
X415 1 3 DCAPBWP7T $T=512280 445080 0 0 $X=511990 $Y=444845
X416 1 3 DCAPBWP7T $T=517880 437240 1 0 $X=517590 $Y=433030
X417 1 3 DCAPBWP7T $T=517880 476440 1 0 $X=517590 $Y=472230
X418 1 3 DCAPBWP7T $T=519000 421560 1 0 $X=518710 $Y=417350
X419 1 3 DCAPBWP7T $T=523480 366680 1 0 $X=523190 $Y=362470
X420 1 3 DCAPBWP7T $T=534120 374520 1 0 $X=533830 $Y=370310
X421 1 3 DCAPBWP7T $T=534120 460760 0 0 $X=533830 $Y=460525
X422 1 3 DCAPBWP7T $T=540840 421560 1 0 $X=540550 $Y=417350
X423 1 3 DCAPBWP7T $T=540840 452920 0 0 $X=540550 $Y=452685
X424 1 3 DCAPBWP7T $T=545320 445080 0 0 $X=545030 $Y=444845
X425 1 3 DCAPBWP7T $T=546440 398040 0 0 $X=546150 $Y=397805
X426 1 3 DCAPBWP7T $T=556520 437240 0 0 $X=556230 $Y=437005
X427 1 3 DCAPBWP7T $T=557080 398040 1 0 $X=556790 $Y=393830
X428 1 3 DCAPBWP7T $T=580600 429400 1 0 $X=580310 $Y=425190
X429 1 3 DCAPBWP7T $T=580600 445080 0 0 $X=580310 $Y=444845
X430 1 3 DCAPBWP7T $T=585080 382360 0 0 $X=584790 $Y=382125
X431 1 3 DCAPBWP7T $T=586760 398040 1 0 $X=586470 $Y=393830
X432 1 3 DCAPBWP7T $T=590680 382360 0 0 $X=590390 $Y=382125
X433 1 3 DCAPBWP7T $T=596280 374520 1 0 $X=595990 $Y=370310
X434 1 3 DCAPBWP7T $T=597960 476440 1 0 $X=597670 $Y=472230
X435 1 3 DCAPBWP7T $T=601320 382360 0 0 $X=601030 $Y=382125
X436 1 3 DCAPBWP7T $T=603000 405880 1 0 $X=602710 $Y=401670
X437 1 3 DCAPBWP7T $T=603000 445080 0 0 $X=602710 $Y=444845
X438 1 3 DCAPBWP7T $T=618120 445080 1 0 $X=617830 $Y=440870
X439 1 3 DCAPBWP7T $T=622600 366680 0 0 $X=622310 $Y=366445
X440 1 3 DCAPBWP7T $T=631000 468600 0 0 $X=630710 $Y=468365
X441 1 3 DCAPBWP7T $T=648360 468600 1 0 $X=648070 $Y=464390
X442 1 3 DCAPBWP7T $T=670760 484280 1 0 $X=670470 $Y=480070
X443 1 3 DCAPBWP7T $T=673560 429400 1 0 $X=673270 $Y=425190
X444 1 3 DCAPBWP7T $T=680280 366680 0 0 $X=679990 $Y=366445
X445 1 3 DCAPBWP7T $T=716680 452920 0 0 $X=716390 $Y=452685
X446 1 3 DCAPBWP7T $T=717800 390200 0 0 $X=717510 $Y=389965
X447 1 3 DCAPBWP7T $T=733480 460760 1 0 $X=733190 $Y=456550
X448 1 3 DCAPBWP7T $T=741320 460760 0 0 $X=741030 $Y=460525
X449 1 3 DCAPBWP7T $T=741320 468600 0 0 $X=741030 $Y=468365
X450 1 3 DCAPBWP7T $T=741320 476440 1 0 $X=741030 $Y=472230
X451 3 1 DCAP8BWP7T $T=458520 445080 1 0 $X=458230 $Y=440870
X452 3 1 DCAP8BWP7T $T=462440 437240 1 0 $X=462150 $Y=433030
X453 3 1 DCAP8BWP7T $T=463560 405880 1 0 $X=463270 $Y=401670
X454 3 1 DCAP8BWP7T $T=464120 390200 1 0 $X=463830 $Y=385990
X455 3 1 DCAP8BWP7T $T=471400 429400 1 0 $X=471110 $Y=425190
X456 3 1 DCAP8BWP7T $T=485960 405880 1 0 $X=485670 $Y=401670
X457 3 1 DCAP8BWP7T $T=485960 421560 0 0 $X=485670 $Y=421325
X458 3 1 DCAP8BWP7T $T=492120 405880 0 0 $X=491830 $Y=405645
X459 3 1 DCAP8BWP7T $T=492120 460760 1 0 $X=491830 $Y=456550
X460 3 1 DCAP8BWP7T $T=494920 445080 0 0 $X=494630 $Y=444845
X461 3 1 DCAP8BWP7T $T=495480 460760 0 0 $X=495190 $Y=460525
X462 3 1 DCAP8BWP7T $T=513400 476440 1 0 $X=513110 $Y=472230
X463 3 1 DCAP8BWP7T $T=526840 476440 1 0 $X=526550 $Y=472230
X464 3 1 DCAP8BWP7T $T=527400 421560 1 0 $X=527110 $Y=417350
X465 3 1 DCAP8BWP7T $T=534120 484280 1 0 $X=533830 $Y=480070
X466 3 1 DCAP8BWP7T $T=546440 460760 0 0 $X=546150 $Y=460525
X467 3 1 DCAP8BWP7T $T=552040 437240 0 0 $X=551750 $Y=437005
X468 3 1 DCAP8BWP7T $T=552040 476440 1 0 $X=551750 $Y=472230
X469 3 1 DCAP8BWP7T $T=562120 445080 0 0 $X=561830 $Y=444845
X470 3 1 DCAP8BWP7T $T=569400 358840 0 0 $X=569110 $Y=358605
X471 3 1 DCAP8BWP7T $T=569400 374520 0 0 $X=569110 $Y=374285
X472 3 1 DCAP8BWP7T $T=569960 405880 0 0 $X=569670 $Y=405645
X473 3 1 DCAP8BWP7T $T=576120 382360 0 0 $X=575830 $Y=382125
X474 3 1 DCAP8BWP7T $T=576120 429400 1 0 $X=575830 $Y=425190
X475 3 1 DCAP8BWP7T $T=576120 437240 0 0 $X=575830 $Y=437005
X476 3 1 DCAP8BWP7T $T=576120 445080 0 0 $X=575830 $Y=444845
X477 3 1 DCAP8BWP7T $T=592920 382360 1 0 $X=592630 $Y=378150
X478 3 1 DCAP8BWP7T $T=593480 476440 1 0 $X=593190 $Y=472230
X479 3 1 DCAP8BWP7T $T=594040 460760 1 0 $X=593750 $Y=456550
X480 3 1 DCAP8BWP7T $T=594600 398040 1 0 $X=594310 $Y=393830
X481 3 1 DCAP8BWP7T $T=601320 382360 1 0 $X=601030 $Y=378150
X482 3 1 DCAP8BWP7T $T=611400 398040 1 0 $X=611110 $Y=393830
X483 3 1 DCAP8BWP7T $T=611400 405880 0 0 $X=611110 $Y=405645
X484 3 1 DCAP8BWP7T $T=611400 445080 0 0 $X=611110 $Y=444845
X485 3 1 DCAP8BWP7T $T=611960 374520 1 0 $X=611670 $Y=370310
X486 3 1 DCAP8BWP7T $T=611960 413720 1 0 $X=611670 $Y=409510
X487 3 1 DCAP8BWP7T $T=611960 468600 1 0 $X=611670 $Y=464390
X488 3 1 DCAP8BWP7T $T=611960 484280 1 0 $X=611670 $Y=480070
X489 3 1 DCAP8BWP7T $T=618120 366680 0 0 $X=617830 $Y=366445
X490 3 1 DCAP8BWP7T $T=618120 429400 0 0 $X=617830 $Y=429165
X491 3 1 DCAP8BWP7T $T=618120 437240 1 0 $X=617830 $Y=433030
X492 3 1 DCAP8BWP7T $T=627080 452920 0 0 $X=626790 $Y=452685
X493 3 1 DCAP8BWP7T $T=639960 445080 1 0 $X=639670 $Y=440870
X494 3 1 DCAP8BWP7T $T=641080 366680 0 0 $X=640790 $Y=366445
X495 3 1 DCAP8BWP7T $T=642760 484280 1 0 $X=642470 $Y=480070
X496 3 1 DCAP8BWP7T $T=643880 468600 1 0 $X=643590 $Y=464390
X497 3 1 DCAP8BWP7T $T=652840 366680 0 0 $X=652550 $Y=366445
X498 3 1 DCAP8BWP7T $T=652840 374520 0 0 $X=652550 $Y=374285
X499 3 1 DCAP8BWP7T $T=653960 374520 1 0 $X=653670 $Y=370310
X500 3 1 DCAP8BWP7T $T=653960 429400 0 0 $X=653670 $Y=429165
X501 3 1 DCAP8BWP7T $T=660120 382360 1 0 $X=659830 $Y=378150
X502 3 1 DCAP8BWP7T $T=660120 437240 1 0 $X=659830 $Y=433030
X503 3 1 DCAP8BWP7T $T=660120 468600 0 0 $X=659830 $Y=468365
X504 3 1 DCAP8BWP7T $T=675800 366680 0 0 $X=675510 $Y=366445
X505 3 1 DCAP8BWP7T $T=694840 366680 1 0 $X=694550 $Y=362470
X506 3 1 DCAP8BWP7T $T=694840 413720 0 0 $X=694550 $Y=413485
X507 3 1 DCAP8BWP7T $T=694840 437240 1 0 $X=694550 $Y=433030
X508 3 1 DCAP8BWP7T $T=695400 445080 1 0 $X=695110 $Y=440870
X509 3 1 DCAP8BWP7T $T=695960 460760 0 0 $X=695670 $Y=460525
X510 3 1 DCAP8BWP7T $T=702120 468600 1 0 $X=701830 $Y=464390
X511 3 1 DCAP8BWP7T $T=706040 413720 1 0 $X=705750 $Y=409510
X512 3 1 DCAP8BWP7T $T=713880 413720 1 0 $X=713590 $Y=409510
X513 3 1 DCAP8BWP7T $T=719480 468600 0 0 $X=719190 $Y=468365
X514 3 1 DCAP8BWP7T $T=723400 413720 1 0 $X=723110 $Y=409510
X515 3 1 DCAP8BWP7T $T=723400 421560 0 0 $X=723110 $Y=421325
X516 3 1 DCAP8BWP7T $T=723400 476440 0 0 $X=723110 $Y=476205
X517 3 1 DCAP8BWP7T $T=736840 468600 0 0 $X=736550 $Y=468365
X518 3 1 DCAP8BWP7T $T=737400 398040 0 0 $X=737110 $Y=397805
X519 3 1 DCAP8BWP7T $T=737960 421560 1 0 $X=737670 $Y=417350
X520 3 1 DCAP8BWP7T $T=737960 429400 1 0 $X=737670 $Y=425190
X521 3 1 DCAP4BWP7T $T=468040 382360 1 0 $X=467750 $Y=378150
X522 3 1 DCAP4BWP7T $T=468040 421560 1 0 $X=467750 $Y=417350
X523 3 1 DCAP4BWP7T $T=488760 460760 1 0 $X=488470 $Y=456550
X524 3 1 DCAP4BWP7T $T=534120 413720 0 0 $X=533830 $Y=413485
X525 3 1 DCAP4BWP7T $T=545320 476440 0 0 $X=545030 $Y=476205
X526 3 1 DCAP4BWP7T $T=557640 413720 1 0 $X=557350 $Y=409510
X527 3 1 DCAP4BWP7T $T=563800 460760 0 0 $X=563510 $Y=460525
X528 3 1 DCAP4BWP7T $T=589560 476440 1 0 $X=589270 $Y=472230
X529 3 1 DCAP4BWP7T $T=618120 405880 1 0 $X=617830 $Y=401670
X530 3 1 DCAP4BWP7T $T=636040 382360 1 0 $X=635750 $Y=378150
X531 3 1 DCAP4BWP7T $T=642760 437240 0 0 $X=642470 $Y=437005
X532 3 1 DCAP4BWP7T $T=645560 429400 0 0 $X=645270 $Y=429165
X533 3 1 DCAP4BWP7T $T=656760 405880 0 0 $X=656470 $Y=405645
X534 3 1 DCAP4BWP7T $T=656760 452920 1 0 $X=656470 $Y=448710
X535 3 1 DCAP4BWP7T $T=660120 398040 1 0 $X=659830 $Y=393830
X536 3 1 DCAP4BWP7T $T=702120 366680 1 0 $X=701830 $Y=362470
X537 3 1 DCAP4BWP7T $T=702120 429400 1 0 $X=701830 $Y=425190
X538 3 1 DCAP4BWP7T $T=740200 390200 0 0 $X=739910 $Y=389965
X539 3 1 DCAP4BWP7T $T=740760 358840 0 0 $X=740470 $Y=358605
X540 3 1 ICV_40 $T=450120 421560 0 0 $X=449830 $Y=421325
X541 3 1 ICV_40 $T=463000 366680 0 0 $X=462710 $Y=366445
X542 3 1 ICV_40 $T=468040 405880 0 0 $X=467750 $Y=405645
X543 3 1 ICV_40 $T=473640 390200 1 0 $X=473350 $Y=385990
X544 3 1 ICV_40 $T=483160 374520 1 0 $X=482870 $Y=370310
X545 3 1 ICV_40 $T=483720 390200 1 0 $X=483430 $Y=385990
X546 3 1 ICV_40 $T=483720 460760 0 0 $X=483430 $Y=460525
X547 3 1 ICV_40 $T=484280 484280 1 0 $X=483990 $Y=480070
X548 3 1 ICV_40 $T=492120 374520 1 0 $X=491830 $Y=370310
X549 3 1 ICV_40 $T=492120 413720 0 0 $X=491830 $Y=413485
X550 3 1 ICV_40 $T=492120 445080 1 0 $X=491830 $Y=440870
X551 3 1 ICV_40 $T=492120 452920 1 0 $X=491830 $Y=448710
X552 3 1 ICV_40 $T=502200 374520 1 0 $X=501910 $Y=370310
X553 3 1 ICV_40 $T=508360 460760 0 0 $X=508070 $Y=460525
X554 3 1 ICV_40 $T=513960 374520 1 0 $X=513670 $Y=370310
X555 3 1 ICV_40 $T=516760 366680 1 0 $X=516470 $Y=362470
X556 3 1 ICV_40 $T=525160 358840 0 0 $X=524870 $Y=358605
X557 3 1 ICV_40 $T=525160 374520 1 0 $X=524870 $Y=370310
X558 3 1 ICV_40 $T=525160 390200 0 0 $X=524870 $Y=389965
X559 3 1 ICV_40 $T=525160 445080 0 0 $X=524870 $Y=444845
X560 3 1 ICV_40 $T=525160 452920 0 0 $X=524870 $Y=452685
X561 3 1 ICV_40 $T=525720 405880 0 0 $X=525430 $Y=405645
X562 3 1 ICV_40 $T=534120 421560 1 0 $X=533830 $Y=417350
X563 3 1 ICV_40 $T=534120 429400 1 0 $X=533830 $Y=425190
X564 3 1 ICV_40 $T=534120 452920 0 0 $X=533830 $Y=452685
X565 3 1 ICV_40 $T=538600 445080 0 0 $X=538310 $Y=444845
X566 3 1 ICV_40 $T=545320 421560 0 0 $X=545030 $Y=421325
X567 3 1 ICV_40 $T=547000 382360 0 0 $X=546710 $Y=382125
X568 3 1 ICV_40 $T=548680 445080 0 0 $X=548390 $Y=444845
X569 3 1 ICV_40 $T=561000 460760 1 0 $X=560710 $Y=456550
X570 3 1 ICV_40 $T=566600 413720 1 0 $X=566310 $Y=409510
X571 3 1 ICV_40 $T=566600 437240 0 0 $X=566310 $Y=437005
X572 3 1 ICV_40 $T=567720 398040 0 0 $X=567430 $Y=397805
X573 3 1 ICV_40 $T=576120 421560 0 0 $X=575830 $Y=421325
X574 3 1 ICV_40 $T=580040 398040 1 0 $X=579750 $Y=393830
X575 3 1 ICV_40 $T=592360 405880 0 0 $X=592070 $Y=405645
X576 3 1 ICV_40 $T=594040 413720 1 0 $X=593750 $Y=409510
X577 3 1 ICV_40 $T=609160 445080 1 0 $X=608870 $Y=440870
X578 3 1 ICV_40 $T=610280 429400 0 0 $X=609990 $Y=429165
X579 3 1 ICV_40 $T=618120 413720 1 0 $X=617830 $Y=409510
X580 3 1 ICV_40 $T=629320 366680 0 0 $X=629030 $Y=366445
X581 3 1 ICV_40 $T=631560 484280 1 0 $X=631270 $Y=480070
X582 3 1 ICV_40 $T=636040 445080 0 0 $X=635750 $Y=444845
X583 3 1 ICV_40 $T=642200 429400 1 0 $X=641910 $Y=425190
X584 3 1 ICV_40 $T=650600 358840 0 0 $X=650310 $Y=358605
X585 3 1 ICV_40 $T=651160 429400 1 0 $X=650870 $Y=425190
X586 3 1 ICV_40 $T=651720 437240 1 0 $X=651430 $Y=433030
X587 3 1 ICV_40 $T=651720 460760 0 0 $X=651430 $Y=460525
X588 3 1 ICV_40 $T=652280 421560 1 0 $X=651990 $Y=417350
X589 3 1 ICV_40 $T=652280 476440 1 0 $X=651990 $Y=472230
X590 3 1 ICV_40 $T=652280 484280 1 0 $X=651990 $Y=480070
X591 3 1 ICV_40 $T=660120 460760 1 0 $X=659830 $Y=456550
X592 3 1 ICV_40 $T=664040 484280 1 0 $X=663750 $Y=480070
X593 3 1 ICV_40 $T=678040 398040 0 0 $X=677750 $Y=397805
X594 3 1 ICV_40 $T=692600 405880 1 0 $X=692310 $Y=401670
X595 3 1 ICV_40 $T=693160 382360 1 0 $X=692870 $Y=378150
X596 3 1 ICV_40 $T=693160 452920 0 0 $X=692870 $Y=452685
X597 3 1 ICV_40 $T=694280 468600 1 0 $X=693990 $Y=464390
X598 3 1 ICV_40 $T=706040 452920 1 0 $X=705750 $Y=448710
X599 3 1 ICV_40 $T=727880 374520 0 0 $X=727590 $Y=374285
X600 3 1 ICV_40 $T=735720 413720 0 0 $X=735430 $Y=413485
X601 21 1 5 8 3 NR2D1BWP7T $T=452920 452920 1 180 $X=450390 $Y=452685
X602 8 1 16 9 3 NR2D1BWP7T $T=452920 460760 0 180 $X=450390 $Y=456550
X603 17 1 22 27 3 NR2D1BWP7T $T=451240 484280 1 0 $X=450950 $Y=480070
X604 42 1 43 27 3 NR2D1BWP7T $T=455720 484280 1 0 $X=455430 $Y=480070
X605 76 1 75 27 3 NR2D1BWP7T $T=484280 484280 0 180 $X=481750 $Y=480070
X606 77 1 78 291 3 NR2D1BWP7T $T=484280 468600 1 0 $X=483990 $Y=464390
X607 294 1 270 27 3 NR2D1BWP7T $T=494920 445080 1 180 $X=492390 $Y=444845
X608 80 1 79 291 3 NR2D1BWP7T $T=495480 460760 1 180 $X=492950 $Y=460525
X609 297 1 285 27 3 NR2D1BWP7T $T=496600 452920 1 180 $X=494070 $Y=452685
X610 291 1 267 27 3 NR2D1BWP7T $T=499960 468600 0 180 $X=497430 $Y=464390
X611 86 1 83 27 3 NR2D1BWP7T $T=500520 468600 1 180 $X=497990 $Y=468365
X612 98 1 286 27 3 NR2D1BWP7T $T=518440 460760 1 180 $X=515910 $Y=460525
X613 332 1 279 27 3 NR2D1BWP7T $T=519000 460760 0 180 $X=516470 $Y=456550
X614 80 1 110 98 3 NR2D1BWP7T $T=524040 460760 0 0 $X=523750 $Y=460525
X615 80 1 340 332 3 NR2D1BWP7T $T=526280 460760 0 0 $X=525990 $Y=460525
X616 112 1 343 291 3 NR2D1BWP7T $T=536920 468600 1 180 $X=534390 $Y=468365
X617 291 1 356 113 3 NR2D1BWP7T $T=539720 484280 1 0 $X=539430 $Y=480070
X618 113 1 115 76 3 NR2D1BWP7T $T=541960 468600 0 0 $X=541670 $Y=468365
X619 86 1 116 113 3 NR2D1BWP7T $T=543080 468600 1 0 $X=542790 $Y=464390
X620 291 1 363 140 3 NR2D1BWP7T $T=545320 468600 1 0 $X=545030 $Y=464390
X621 113 1 364 98 3 NR2D1BWP7T $T=546440 452920 1 0 $X=546150 $Y=448710
X622 358 1 383 368 3 NR2D1BWP7T $T=560440 437240 1 0 $X=560150 $Y=433030
X623 86 1 380 135 3 NR2D1BWP7T $T=566040 460760 0 0 $X=565750 $Y=460525
X624 297 1 373 77 3 NR2D1BWP7T $T=570520 452920 0 180 $X=567990 $Y=448710
X625 80 1 399 297 3 NR2D1BWP7T $T=568280 460760 1 0 $X=567990 $Y=456550
X626 77 1 388 332 3 NR2D1BWP7T $T=568280 460760 0 0 $X=567990 $Y=460525
X627 86 1 365 140 3 NR2D1BWP7T $T=578920 452920 1 0 $X=578630 $Y=448710
X628 130 1 419 133 3 NR2D1BWP7T $T=581720 382360 1 0 $X=581430 $Y=378150
X629 112 1 412 98 3 NR2D1BWP7T $T=581720 452920 1 0 $X=581430 $Y=448710
X630 80 1 384 294 3 NR2D1BWP7T $T=583960 452920 1 0 $X=583670 $Y=448710
X631 112 1 422 332 3 NR2D1BWP7T $T=585080 445080 0 0 $X=584790 $Y=444845
X632 1 3 DCAP64BWP7T $T=452920 460760 1 0 $X=452630 $Y=456550
X633 1 3 DCAP64BWP7T $T=453480 452920 1 0 $X=453190 $Y=448710
X634 1 3 DCAP64BWP7T $T=538040 429400 0 0 $X=537750 $Y=429165
X635 1 3 DCAP64BWP7T $T=539160 413720 0 0 $X=538870 $Y=413485
X684 3 1 ICV_47 $T=450120 390200 0 0 $X=449830 $Y=389965
X685 3 1 ICV_47 $T=450120 429400 0 0 $X=449830 $Y=429165
X686 3 1 ICV_47 $T=492120 429400 1 0 $X=491830 $Y=425190
X687 3 1 ICV_47 $T=492120 429400 0 0 $X=491830 $Y=429165
X688 3 1 ICV_47 $T=492120 437240 0 0 $X=491830 $Y=437005
X689 3 1 ICV_47 $T=534120 390200 0 0 $X=533830 $Y=389965
X690 3 1 ICV_47 $T=534120 405880 1 0 $X=533830 $Y=401670
X691 3 1 ICV_47 $T=534120 445080 1 0 $X=533830 $Y=440870
X692 3 1 ICV_47 $T=576120 366680 1 0 $X=575830 $Y=362470
X693 3 1 ICV_47 $T=576120 468600 0 0 $X=575830 $Y=468365
X694 3 1 ICV_47 $T=576120 476440 0 0 $X=575830 $Y=476205
X695 3 1 ICV_47 $T=618120 382360 0 0 $X=617830 $Y=382125
X696 3 1 ICV_47 $T=618120 398040 0 0 $X=617830 $Y=397805
X697 3 1 ICV_47 $T=660120 429400 0 0 $X=659830 $Y=429165
X698 3 1 ICV_47 $T=660120 476440 0 0 $X=659830 $Y=476205
X699 3 1 ICV_47 $T=702120 484280 1 0 $X=701830 $Y=480070
X700 1 3 DCAP32BWP7T $T=450120 382360 1 0 $X=449830 $Y=378150
X701 1 3 DCAP32BWP7T $T=450120 405880 0 0 $X=449830 $Y=405645
X702 1 3 DCAP32BWP7T $T=450120 421560 1 0 $X=449830 $Y=417350
X703 1 3 DCAP32BWP7T $T=450120 460760 0 0 $X=449830 $Y=460525
X704 1 3 DCAP32BWP7T $T=458520 366680 1 0 $X=458230 $Y=362470
X705 1 3 DCAP32BWP7T $T=461880 398040 0 0 $X=461590 $Y=397805
X706 1 3 DCAP32BWP7T $T=465240 374520 1 0 $X=464950 $Y=370310
X707 1 3 DCAP32BWP7T $T=468040 421560 0 0 $X=467750 $Y=421325
X708 1 3 DCAP32BWP7T $T=492120 413720 1 0 $X=491830 $Y=409510
X709 1 3 DCAP32BWP7T $T=503320 445080 1 0 $X=503030 $Y=440870
X710 1 3 DCAP32BWP7T $T=507240 452920 0 0 $X=506950 $Y=452685
X711 1 3 DCAP32BWP7T $T=534120 358840 0 0 $X=533830 $Y=358605
X712 1 3 DCAP32BWP7T $T=534120 398040 1 0 $X=533830 $Y=393830
X713 1 3 DCAP32BWP7T $T=534120 476440 1 0 $X=533830 $Y=472230
X714 1 3 DCAP32BWP7T $T=551480 374520 0 0 $X=551190 $Y=374285
X715 1 3 DCAP32BWP7T $T=557080 421560 1 0 $X=556790 $Y=417350
X716 1 3 DCAP32BWP7T $T=576120 390200 0 0 $X=575830 $Y=389965
X717 1 3 DCAP32BWP7T $T=576120 413720 1 0 $X=575830 $Y=409510
X718 1 3 DCAP32BWP7T $T=576120 429400 0 0 $X=575830 $Y=429165
X719 1 3 DCAP32BWP7T $T=576120 460760 1 0 $X=575830 $Y=456550
X720 1 3 DCAP32BWP7T $T=618120 358840 0 0 $X=617830 $Y=358605
X721 1 3 DCAP32BWP7T $T=618120 445080 0 0 $X=617830 $Y=444845
X722 1 3 DCAP32BWP7T $T=618120 476440 0 0 $X=617830 $Y=476205
X723 1 3 DCAP32BWP7T $T=624280 429400 1 0 $X=623990 $Y=425190
X724 1 3 DCAP32BWP7T $T=634360 421560 1 0 $X=634070 $Y=417350
X725 1 3 DCAP32BWP7T $T=636040 374520 1 0 $X=635750 $Y=370310
X726 1 3 DCAP32BWP7T $T=639960 476440 0 0 $X=639670 $Y=476205
X727 1 3 DCAP32BWP7T $T=660120 366680 1 0 $X=659830 $Y=362470
X728 1 3 DCAP32BWP7T $T=660120 374520 1 0 $X=659830 $Y=370310
X729 1 3 DCAP32BWP7T $T=660120 398040 0 0 $X=659830 $Y=397805
X730 1 3 DCAP32BWP7T $T=660120 452920 1 0 $X=659830 $Y=448710
X731 1 3 DCAP32BWP7T $T=671880 405880 0 0 $X=671590 $Y=405645
X732 1 3 DCAP32BWP7T $T=675240 382360 1 0 $X=674950 $Y=378150
X733 1 3 DCAP32BWP7T $T=675240 452920 0 0 $X=674950 $Y=452685
X734 1 3 DCAP32BWP7T $T=676360 468600 1 0 $X=676070 $Y=464390
X735 1 3 DCAP32BWP7T $T=702120 405880 0 0 $X=701830 $Y=405645
X736 1 3 DCAP32BWP7T $T=702120 421560 1 0 $X=701830 $Y=417350
X737 1 3 DCAP32BWP7T $T=702120 437240 1 0 $X=701830 $Y=433030
X738 1 3 DCAP32BWP7T $T=702120 445080 0 0 $X=701830 $Y=444845
X739 1 3 DCAP32BWP7T $T=702120 460760 1 0 $X=701830 $Y=456550
X740 1 3 DCAP32BWP7T $T=719480 398040 0 0 $X=719190 $Y=397805
X741 1 3 DCAP32BWP7T $T=722280 390200 0 0 $X=721990 $Y=389965
X742 1 3 DCAP32BWP7T $T=722840 358840 0 0 $X=722550 $Y=358605
X743 10 37 47 55 1 3 56 FA1D0BWP7T $T=450680 468600 1 0 $X=450390 $Y=464390
X744 365 343 340 129 1 3 132 FA1D0BWP7T $T=547560 476440 0 0 $X=547270 $Y=476205
X745 373 126 384 390 1 3 393 FA1D0BWP7T $T=550920 460760 0 0 $X=550630 $Y=460525
X746 380 388 399 137 1 3 405 FA1D0BWP7T $T=557640 476440 1 0 $X=557350 $Y=472230
X747 138 412 356 148 1 3 428 FA1D0BWP7T $T=576680 476440 1 0 $X=576390 $Y=472230
X748 364 363 422 427 1 3 429 FA1D0BWP7T $T=577240 460760 0 0 $X=576950 $Y=460525
X749 390 428 427 435 1 3 438 FA1D0BWP7T $T=590120 468600 1 0 $X=589830 $Y=464390
X750 152 405 154 436 1 3 443 FA1D0BWP7T $T=590120 484280 1 0 $X=589830 $Y=480070
X751 435 436 164 163 1 3 448 FA1D0BWP7T $T=631560 484280 0 180 $X=618390 $Y=480070
X752 102 3 1 291 INVD1BWP7T $T=593480 476440 0 180 $X=591510 $Y=472230
X753 124 3 1 156 INVD1BWP7T $T=606360 405880 0 180 $X=604390 $Y=401670
X754 172 3 1 98 INVD1BWP7T $T=633240 452920 1 180 $X=631270 $Y=452685
X755 198 3 1 297 INVD1BWP7T $T=651160 429400 0 180 $X=649190 $Y=425190
X756 452 3 1 186 CKBD0BWP7T $T=641640 468600 1 0 $X=641350 $Y=464390
X875 24 3 20 15 1 ND2D1BWP7T $T=453480 452920 0 180 $X=450950 $Y=448710
X876 36 3 30 23 1 ND2D1BWP7T $T=455160 445080 0 180 $X=452630 $Y=440870
X877 32 3 35 246 1 ND2D1BWP7T $T=453480 484280 1 0 $X=453190 $Y=480070
X878 51 3 255 256 1 ND2D1BWP7T $T=461320 437240 0 0 $X=461030 $Y=437005
X879 66 3 262 64 1 ND2D1BWP7T $T=470840 437240 0 180 $X=468310 $Y=433030
X880 65 3 73 85 1 ND2D1BWP7T $T=497720 460760 1 0 $X=497430 $Y=456550
X881 316 3 87 273 1 ND2D1BWP7T $T=508360 460760 1 180 $X=505830 $Y=460525
X882 100 3 104 108 1 ND2D1BWP7T $T=522360 476440 1 0 $X=522070 $Y=472230
X883 100 3 105 111 1 ND2D1BWP7T $T=522360 484280 1 0 $X=522070 $Y=480070
X884 303 3 351 369 1 ND2D1BWP7T $T=552040 437240 1 180 $X=549510 $Y=437005
X885 342 3 358 345 1 ND2D1BWP7T $T=559880 445080 0 0 $X=559590 $Y=444845
X886 131 3 396 100 1 ND2D1BWP7T $T=566600 437240 1 180 $X=564070 $Y=437005
X887 85 3 381 352 1 ND2D1BWP7T $T=577240 413720 0 0 $X=576950 $Y=413485
X888 441 3 406 430 1 ND2D1BWP7T $T=605240 382360 1 180 $X=602710 $Y=382125
X889 133 3 440 130 1 ND2D1BWP7T $T=620920 390200 0 180 $X=618390 $Y=385990
X890 162 3 449 161 1 ND2D1BWP7T $T=623720 445080 0 180 $X=621190 $Y=440870
X891 142 3 431 111 1 ND2D1BWP7T $T=624840 437240 0 180 $X=622310 $Y=433030
X892 102 3 444 167 1 ND2D1BWP7T $T=622600 460760 0 0 $X=622310 $Y=460525
X893 174 3 447 172 1 ND2D1BWP7T $T=633800 460760 0 180 $X=631270 $Y=456550
X894 211 3 516 212 1 ND2D1BWP7T $T=678040 382360 0 0 $X=677750 $Y=382125
X895 211 3 220 221 1 ND2D1BWP7T $T=702680 366680 0 0 $X=702390 $Y=366445
X923 246 3 1 42 INVD0BWP7T $T=458520 445080 0 180 $X=456550 $Y=440870
X924 67 3 1 68 INVD0BWP7T $T=470280 468600 1 0 $X=469990 $Y=464390
X925 273 3 1 271 INVD0BWP7T $T=477000 452920 1 180 $X=475030 $Y=452685
X926 292 3 1 293 INVD0BWP7T $T=492680 452920 0 0 $X=492390 $Y=452685
X927 87 3 1 321 INVD0BWP7T $T=515640 468600 1 180 $X=513670 $Y=468365
X928 314 3 1 359 INVD0BWP7T $T=534680 421560 0 0 $X=534390 $Y=421325
X929 361 3 1 360 INVD0BWP7T $T=547000 382360 1 180 $X=545030 $Y=382125
X930 344 3 1 348 INVD0BWP7T $T=547560 437240 0 180 $X=545590 $Y=433030
X931 367 3 1 368 INVD0BWP7T $T=548680 437240 1 0 $X=548390 $Y=433030
X932 376 3 1 378 INVD0BWP7T $T=557080 398040 0 180 $X=555110 $Y=393830
X933 397 3 1 395 INVD0BWP7T $T=567160 382360 1 180 $X=565190 $Y=382125
X934 394 3 1 401 INVD0BWP7T $T=576680 437240 1 0 $X=576390 $Y=433030
X935 433 3 1 413 INVD0BWP7T $T=606920 421560 0 180 $X=604950 $Y=417350
X936 162 3 1 294 INVD0BWP7T $T=611400 445080 1 180 $X=609430 $Y=444845
X937 6 13 18 25 3 1 OAI21D0BWP7T $T=450680 374520 1 0 $X=450390 $Y=370310
X938 26 244 18 7 3 1 OAI21D0BWP7T $T=453480 382360 1 180 $X=450390 $Y=382125
X939 39 250 48 253 3 1 OAI21D0BWP7T $T=459080 413720 0 0 $X=458790 $Y=413485
X940 45 251 18 248 3 1 OAI21D0BWP7T $T=463000 366680 1 180 $X=459910 $Y=366445
X941 48 252 53 258 3 1 OAI21D0BWP7T $T=460760 405880 1 0 $X=460470 $Y=401670
X942 26 260 48 259 3 1 OAI21D0BWP7T $T=461320 382360 0 0 $X=461030 $Y=382125
X943 6 247 48 261 3 1 OAI21D0BWP7T $T=462440 374520 1 0 $X=462150 $Y=370310
X944 39 249 70 274 3 1 OAI21D0BWP7T $T=474200 413720 1 0 $X=473910 $Y=409510
X945 70 266 53 276 3 1 OAI21D0BWP7T $T=475880 405880 0 0 $X=475590 $Y=405645
X946 48 278 72 280 3 1 OAI21D0BWP7T $T=486520 358840 1 180 $X=483430 $Y=358605
X947 45 283 48 264 3 1 OAI21D0BWP7T $T=486520 366680 1 180 $X=483430 $Y=366445
X948 26 287 70 281 3 1 OAI21D0BWP7T $T=496040 398040 0 180 $X=492950 $Y=393830
X949 39 296 81 289 3 1 OAI21D0BWP7T $T=496600 405880 0 180 $X=493510 $Y=401670
X950 6 295 70 300 3 1 OAI21D0BWP7T $T=495480 374520 0 0 $X=495190 $Y=374285
X951 45 82 70 84 3 1 OAI21D0BWP7T $T=496040 366680 1 0 $X=495750 $Y=362470
X952 81 299 53 301 3 1 OAI21D0BWP7T $T=497160 398040 0 0 $X=496870 $Y=397805
X953 39 304 88 298 3 1 OAI21D0BWP7T $T=502760 413720 1 180 $X=499670 $Y=413485
X954 292 302 303 306 3 1 OAI21D0BWP7T $T=500520 452920 1 0 $X=500230 $Y=448710
X955 26 318 81 308 3 1 OAI21D0BWP7T $T=501080 390200 0 0 $X=500790 $Y=389965
X956 6 313 81 317 3 1 OAI21D0BWP7T $T=506120 382360 1 0 $X=505830 $Y=378150
X957 88 326 53 320 3 1 OAI21D0BWP7T $T=514520 413720 0 180 $X=511430 $Y=409510
X958 45 322 88 106 3 1 OAI21D0BWP7T $T=513400 358840 0 0 $X=513110 $Y=358605
X959 275 324 316 95 3 1 OAI21D0BWP7T $T=516200 460760 0 180 $X=513110 $Y=456550
X960 6 338 88 334 3 1 OAI21D0BWP7T $T=528520 382360 0 180 $X=525430 $Y=378150
X961 26 339 88 336 3 1 OAI21D0BWP7T $T=528520 398040 0 180 $X=525430 $Y=393830
X962 45 346 81 337 3 1 OAI21D0BWP7T $T=537480 366680 0 180 $X=534390 $Y=362470
X963 297 404 112 396 3 1 OAI21D0BWP7T $T=585080 445080 1 180 $X=581990 $Y=444845
X964 433 434 417 421 3 1 OAI21D0BWP7T $T=605240 421560 0 180 $X=602150 $Y=417350
X965 332 451 113 449 3 1 OAI21D0BWP7T $T=622040 452920 0 0 $X=621750 $Y=452685
X966 182 487 184 474 3 1 OAI21D0BWP7T $T=641080 452920 0 0 $X=640790 $Y=452685
X967 191 489 184 478 3 1 OAI21D0BWP7T $T=652840 366680 1 180 $X=649750 $Y=366445
X968 182 490 200 486 3 1 OAI21D0BWP7T $T=652840 468600 0 180 $X=649750 $Y=464390
X969 184 492 482 485 3 1 OAI21D0BWP7T $T=653960 429400 1 180 $X=650870 $Y=429165
X970 188 205 194 206 3 1 OAI21D0BWP7T $T=661240 484280 1 0 $X=660950 $Y=480070
X971 200 497 482 496 3 1 OAI21D0BWP7T $T=661800 452920 0 0 $X=661510 $Y=452685
X972 193 499 184 477 3 1 OAI21D0BWP7T $T=666840 382360 1 180 $X=663750 $Y=382125
X973 483 500 184 493 3 1 OAI21D0BWP7T $T=666840 413720 0 180 $X=663750 $Y=409510
X974 480 501 184 494 3 1 OAI21D0BWP7T $T=666840 421560 0 180 $X=663750 $Y=417350
X975 182 502 207 498 3 1 OAI21D0BWP7T $T=669640 468600 1 180 $X=666550 $Y=468365
X976 193 504 516 506 3 1 OAI21D0BWP7T $T=671880 390200 1 0 $X=671590 $Y=385990
X977 207 503 482 508 3 1 OAI21D0BWP7T $T=672440 452920 0 0 $X=672150 $Y=452685
X978 483 505 200 511 3 1 OAI21D0BWP7T $T=673000 398040 1 0 $X=672710 $Y=393830
X979 480 519 200 507 3 1 OAI21D0BWP7T $T=680840 421560 0 180 $X=677750 $Y=417350
X980 182 213 516 510 3 1 OAI21D0BWP7T $T=681960 468600 1 180 $X=678870 $Y=468365
X981 516 518 191 522 3 1 OAI21D0BWP7T $T=681960 366680 0 0 $X=681670 $Y=366445
X982 480 521 516 528 3 1 OAI21D0BWP7T $T=685320 437240 1 0 $X=685030 $Y=433030
X983 483 523 516 532 3 1 OAI21D0BWP7T $T=688680 429400 1 0 $X=688390 $Y=425190
X984 480 524 207 527 3 1 OAI21D0BWP7T $T=693720 421560 1 180 $X=690630 $Y=421325
X985 182 536 217 537 3 1 OAI21D0BWP7T $T=693160 460760 0 0 $X=692870 $Y=460525
X986 483 535 207 542 3 1 OAI21D0BWP7T $T=693720 390200 0 0 $X=693430 $Y=389965
X987 516 530 482 531 3 1 OAI21D0BWP7T $T=693720 445080 0 0 $X=693430 $Y=444845
X988 480 540 217 553 3 1 OAI21D0BWP7T $T=702680 421560 0 0 $X=702390 $Y=421325
X989 217 541 482 539 3 1 OAI21D0BWP7T $T=703240 452920 1 0 $X=702950 $Y=448710
X990 483 546 217 550 3 1 OAI21D0BWP7T $T=707160 405880 1 0 $X=706870 $Y=401670
X991 182 551 223 552 3 1 OAI21D0BWP7T $T=711640 468600 1 0 $X=711350 $Y=464390
X992 182 222 224 225 3 1 OAI21D0BWP7T $T=711640 476440 1 0 $X=711350 $Y=472230
X993 223 561 482 558 3 1 OAI21D0BWP7T $T=715000 445080 0 180 $X=711910 $Y=440870
X994 223 544 191 563 3 1 OAI21D0BWP7T $T=713320 358840 0 0 $X=713030 $Y=358605
X995 480 549 223 560 3 1 OAI21D0BWP7T $T=716680 429400 1 180 $X=713590 $Y=429165
X996 193 545 220 567 3 1 OAI21D0BWP7T $T=716680 398040 0 0 $X=716390 $Y=397805
X997 224 565 482 568 3 1 OAI21D0BWP7T $T=716680 468600 0 0 $X=716390 $Y=468365
X998 193 572 223 569 3 1 OAI21D0BWP7T $T=722280 390200 1 180 $X=719190 $Y=389965
X999 483 571 223 577 3 1 OAI21D0BWP7T $T=720040 405880 1 0 $X=719750 $Y=401670
X1000 483 548 224 574 3 1 OAI21D0BWP7T $T=720600 413720 1 0 $X=720310 $Y=409510
X1001 480 582 224 579 3 1 OAI21D0BWP7T $T=726200 445080 1 180 $X=723110 $Y=444845
X1002 220 584 482 588 3 1 OAI21D0BWP7T $T=725080 468600 0 0 $X=724790 $Y=468365
X1003 483 590 220 578 3 1 OAI21D0BWP7T $T=737960 421560 0 180 $X=734870 $Y=417350
X1004 220 589 191 559 3 1 OAI21D0BWP7T $T=738520 374520 1 180 $X=735430 $Y=374285
X1005 480 591 220 585 3 1 OAI21D0BWP7T $T=738520 437240 0 180 $X=735430 $Y=433030
X1059 85 3 303 292 1 306 ND3D0BWP7T $T=503320 445080 1 180 $X=500230 $Y=444845
X1060 99 3 100 102 1 103 ND3D0BWP7T $T=519560 476440 1 0 $X=519270 $Y=472230
X1061 3 1 DCAP16BWP7T $T=450120 358840 0 0 $X=449830 $Y=358605
X1062 3 1 DCAP16BWP7T $T=450120 405880 1 0 $X=449830 $Y=401670
X1063 3 1 DCAP16BWP7T $T=450120 413720 0 0 $X=449830 $Y=413485
X1064 3 1 DCAP16BWP7T $T=453480 374520 1 0 $X=453190 $Y=370310
X1065 3 1 DCAP16BWP7T $T=457960 429400 1 0 $X=457670 $Y=425190
X1066 3 1 DCAP16BWP7T $T=468040 484280 1 0 $X=467750 $Y=480070
X1067 3 1 DCAP16BWP7T $T=470280 358840 0 0 $X=469990 $Y=358605
X1068 3 1 DCAP16BWP7T $T=471960 468600 1 0 $X=471670 $Y=464390
X1069 3 1 DCAP16BWP7T $T=473640 405880 1 0 $X=473350 $Y=401670
X1070 3 1 DCAP16BWP7T $T=478680 405880 0 0 $X=478390 $Y=405645
X1071 3 1 DCAP16BWP7T $T=482040 382360 0 0 $X=481750 $Y=382125
X1072 3 1 DCAP16BWP7T $T=492120 366680 0 0 $X=491830 $Y=366445
X1073 3 1 DCAP16BWP7T $T=492120 382360 1 0 $X=491830 $Y=378150
X1074 3 1 DCAP16BWP7T $T=492120 390200 0 0 $X=491830 $Y=389965
X1075 3 1 DCAP16BWP7T $T=500520 468600 0 0 $X=500230 $Y=468365
X1076 3 1 DCAP16BWP7T $T=503320 445080 0 0 $X=503030 $Y=444845
X1077 3 1 DCAP16BWP7T $T=520120 382360 0 0 $X=519830 $Y=382125
X1078 3 1 DCAP16BWP7T $T=534120 374520 0 0 $X=533830 $Y=374285
X1079 3 1 DCAP16BWP7T $T=534120 437240 1 0 $X=533830 $Y=433030
X1080 3 1 DCAP16BWP7T $T=576120 366680 0 0 $X=575830 $Y=366445
X1081 3 1 DCAP16BWP7T $T=576120 468600 1 0 $X=575830 $Y=464390
X1082 3 1 DCAP16BWP7T $T=576120 484280 1 0 $X=575830 $Y=480070
X1083 3 1 DCAP16BWP7T $T=579480 413720 0 0 $X=579190 $Y=413485
X1084 3 1 DCAP16BWP7T $T=603560 358840 0 0 $X=603270 $Y=358605
X1085 3 1 DCAP16BWP7T $T=606360 390200 0 0 $X=606070 $Y=389965
X1086 3 1 DCAP16BWP7T $T=606360 405880 1 0 $X=606070 $Y=401670
X1087 3 1 DCAP16BWP7T $T=618120 374520 1 0 $X=617830 $Y=370310
X1088 3 1 DCAP16BWP7T $T=618120 398040 1 0 $X=617830 $Y=393830
X1089 3 1 DCAP16BWP7T $T=624280 468600 1 0 $X=623990 $Y=464390
X1090 3 1 DCAP16BWP7T $T=634360 366680 1 0 $X=634070 $Y=362470
X1091 3 1 DCAP16BWP7T $T=646120 445080 0 0 $X=645830 $Y=444845
X1092 3 1 DCAP16BWP7T $T=648920 437240 0 0 $X=648630 $Y=437005
X1093 3 1 DCAP16BWP7T $T=648920 468600 0 0 $X=648630 $Y=468365
X1094 3 1 DCAP16BWP7T $T=650040 390200 1 0 $X=649750 $Y=385990
X1095 3 1 DCAP16BWP7T $T=650040 398040 1 0 $X=649750 $Y=393830
X1096 3 1 DCAP16BWP7T $T=669640 468600 0 0 $X=669350 $Y=468365
X1097 3 1 DCAP16BWP7T $T=675240 437240 1 0 $X=674950 $Y=433030
X1098 3 1 DCAP16BWP7T $T=687560 374520 0 0 $X=687270 $Y=374285
X1099 3 1 DCAP16BWP7T $T=690360 421560 1 0 $X=690070 $Y=417350
X1100 3 1 DCAP16BWP7T $T=691480 429400 1 0 $X=691190 $Y=425190
X1101 3 1 DCAP16BWP7T $T=692040 484280 1 0 $X=691750 $Y=480070
X1102 3 1 DCAP16BWP7T $T=702120 374520 0 0 $X=701830 $Y=374285
X1103 3 1 DCAP16BWP7T $T=702120 445080 1 0 $X=701830 $Y=440870
X1104 3 1 DCAP16BWP7T $T=702120 476440 1 0 $X=701830 $Y=472230
X1105 3 1 DCAP16BWP7T $T=706040 460760 0 0 $X=705750 $Y=460525
X1106 3 1 DCAP16BWP7T $T=709960 405880 1 0 $X=709670 $Y=401670
X1107 3 1 DCAP16BWP7T $T=716120 452920 1 0 $X=715830 $Y=448710
X1108 3 1 DCAP16BWP7T $T=718360 437240 0 0 $X=718070 $Y=437005
X1109 3 1 DCAP16BWP7T $T=722840 405880 1 0 $X=722550 $Y=401670
X1110 3 1 DCAP16BWP7T $T=726200 421560 1 0 $X=725910 $Y=417350
X1111 3 1 DCAP16BWP7T $T=729560 429400 0 0 $X=729270 $Y=429165
X1112 3 1 DCAP16BWP7T $T=732920 366680 1 0 $X=732630 $Y=362470
X1113 3 1 DCAP16BWP7T $T=733480 390200 1 0 $X=733190 $Y=385990
X1137 143 3 433 139 394 1 NR3D1BWP7T $T=602440 437240 1 180 $X=597670 $Y=437005
X1138 354 303 3 94 371 1 AOI21D1BWP7T $T=552040 405880 1 180 $X=548390 $Y=405645
X1139 394 402 3 156 158 1 AOI21D1BWP7T $T=608040 445080 1 180 $X=604390 $Y=444845
X1140 245 31 1 3 INVD2BWP7T $T=455160 452920 1 180 $X=452630 $Y=452685
X1141 57 59 1 3 INVD2BWP7T $T=464680 468600 1 0 $X=464390 $Y=464390
X1142 100 80 1 3 INVD2BWP7T $T=523480 460760 1 180 $X=520950 $Y=460525
X1143 108 76 1 3 INVD2BWP7T $T=526840 476440 0 180 $X=524310 $Y=472230
X1144 95 309 1 3 INVD2BWP7T $T=536920 437240 1 180 $X=534390 $Y=437005
X1145 111 86 1 3 INVD2BWP7T $T=535240 452920 1 0 $X=534950 $Y=448710
X1146 327 303 1 3 INVD2BWP7T $T=535800 429400 0 0 $X=535510 $Y=429165
X1147 125 133 1 3 INVD2BWP7T $T=583400 374520 0 0 $X=583110 $Y=374285
X1148 161 77 1 3 INVD2BWP7T $T=609160 445080 0 180 $X=606630 $Y=440870
X1149 446 421 1 3 INVD2BWP7T $T=622040 429400 1 0 $X=621750 $Y=425190
X1150 168 113 1 3 INVD2BWP7T $T=624840 452920 0 0 $X=624550 $Y=452685
X1151 185 332 1 3 INVD2BWP7T $T=643880 374520 1 180 $X=641350 $Y=374285
X1213 34 244 3 1 14 DFQD0BWP7T $T=461880 398040 1 180 $X=450950 $Y=397805
X1214 34 249 3 1 11 DFQD0BWP7T $T=462440 437240 0 180 $X=451510 $Y=433030
X1215 34 251 3 1 28 DFQD0BWP7T $T=464120 374520 1 180 $X=453190 $Y=374285
X1216 34 247 3 1 257 DFQD0BWP7T $T=453480 390200 1 0 $X=453190 $Y=385990
X1217 34 60 3 1 38 DFQD0BWP7T $T=470280 358840 1 180 $X=459350 $Y=358605
X1218 34 252 3 1 263 DFQD0BWP7T $T=459640 413720 1 0 $X=459350 $Y=409510
X1219 34 260 3 1 268 DFQD0BWP7T $T=463560 398040 1 0 $X=463270 $Y=393830
X1220 69 267 3 1 49 DFQD0BWP7T $T=475880 476440 1 180 $X=464950 $Y=476205
X1221 34 266 3 1 282 DFQD0BWP7T $T=470280 421560 1 0 $X=469990 $Y=417350
X1222 34 278 3 1 269 DFQD0BWP7T $T=483720 366680 1 180 $X=472790 $Y=366445
X1223 69 279 3 1 15 DFQD0BWP7T $T=483720 460760 1 180 $X=472790 $Y=460525
X1224 34 283 3 1 265 DFQD0BWP7T $T=486520 382360 0 180 $X=475590 $Y=378150
X1225 34 287 3 1 272 DFQD0BWP7T $T=486520 398040 0 180 $X=475590 $Y=393830
X1226 34 284 3 1 66 DFQD0BWP7T $T=486520 437240 0 180 $X=475590 $Y=433030
X1227 34 285 3 1 36 DFQD0BWP7T $T=486520 445080 1 180 $X=475590 $Y=444845
X1228 69 286 3 1 245 DFQD0BWP7T $T=486520 476440 0 180 $X=475590 $Y=472230
X1229 34 295 3 1 288 DFQD0BWP7T $T=492680 382360 0 0 $X=492390 $Y=382125
X1230 69 277 3 1 273 DFQD0BWP7T $T=493800 476440 1 0 $X=493510 $Y=472230
X1231 34 299 3 1 290 DFQD0BWP7T $T=498280 405880 0 0 $X=497990 $Y=405645
X1232 34 302 3 1 327 DFQD0BWP7T $T=503320 437240 1 0 $X=503030 $Y=433030
X1233 34 313 3 1 323 DFQD0BWP7T $T=505000 382360 0 0 $X=504710 $Y=382125
X1234 34 326 3 1 315 DFQD0BWP7T $T=517880 421560 1 180 $X=506950 $Y=421325
X1235 69 319 3 1 316 DFQD0BWP7T $T=518440 476440 1 180 $X=507510 $Y=476205
X1236 34 318 3 1 328 DFQD0BWP7T $T=508920 398040 1 0 $X=508630 $Y=393830
X1237 34 322 3 1 101 DFQD0BWP7T $T=510600 366680 0 0 $X=510310 $Y=366445
X1238 34 338 3 1 333 DFQD0BWP7T $T=545320 390200 0 180 $X=534390 $Y=385990
X1239 118 357 3 1 342 DFQD0BWP7T $T=545320 476440 1 180 $X=534390 $Y=476205
X1240 34 346 3 1 325 DFQD0BWP7T $T=546440 374520 0 180 $X=535510 $Y=370310
X1241 34 339 3 1 329 DFQD0BWP7T $T=546440 398040 1 180 $X=535510 $Y=397805
X1242 118 349 3 1 344 DFQD0BWP7T $T=546440 460760 1 180 $X=535510 $Y=460525
X1243 34 355 3 1 367 DFQD0BWP7T $T=538600 437240 0 0 $X=538310 $Y=437005
X1244 34 375 3 1 389 DFQD0BWP7T $T=552040 421560 0 0 $X=551750 $Y=421325
X1245 118 387 3 1 369 DFQD0BWP7T $T=564360 452920 0 180 $X=553430 $Y=448710
X1246 118 497 3 1 491 DFQD0BWP7T $T=660680 445080 0 0 $X=660390 $Y=444845
X1247 118 500 3 1 488 DFQD0BWP7T $T=671880 405880 1 180 $X=660950 $Y=405645
X1248 118 501 3 1 481 DFQD0BWP7T $T=672440 421560 1 180 $X=661510 $Y=421325
X1249 118 499 3 1 476 DFQD0BWP7T $T=673000 398040 0 180 $X=662070 $Y=393830
X1250 118 489 3 1 475 DFQD0BWP7T $T=675240 382360 0 180 $X=664310 $Y=378150
X1251 118 492 3 1 479 DFQD0BWP7T $T=675240 437240 0 180 $X=664310 $Y=433030
X1252 118 495 3 1 484 DFQD0BWP7T $T=675800 366680 1 180 $X=664870 $Y=366445
X1253 118 503 3 1 513 DFQD0BWP7T $T=667960 460760 1 0 $X=667670 $Y=456550
X1254 118 505 3 1 514 DFQD0BWP7T $T=673000 405880 1 0 $X=672710 $Y=401670
X1255 118 519 3 1 509 DFQD0BWP7T $T=685880 429400 0 180 $X=674950 $Y=425190
X1256 210 517 3 1 529 DFQD0BWP7T $T=676920 358840 0 0 $X=676630 $Y=358605
X1257 118 518 3 1 526 DFQD0BWP7T $T=676920 374520 0 0 $X=676630 $Y=374285
X1258 118 524 3 1 515 DFQD0BWP7T $T=689240 437240 1 180 $X=678310 $Y=437005
X1259 118 530 3 1 512 DFQD0BWP7T $T=692040 460760 1 180 $X=681110 $Y=460525
X1260 118 521 3 1 533 DFQD0BWP7T $T=681960 452920 1 0 $X=681670 $Y=448710
X1261 118 523 3 1 534 DFQD0BWP7T $T=683080 413720 1 0 $X=682790 $Y=409510
X1262 118 504 3 1 520 DFQD0BWP7T $T=696520 382360 1 180 $X=685590 $Y=382125
X1263 118 535 3 1 525 DFQD0BWP7T $T=696520 398040 1 180 $X=685590 $Y=397805
X1264 210 544 3 1 573 DFQD0BWP7T $T=704360 366680 1 0 $X=704070 $Y=362470
X1265 118 540 3 1 543 DFQD0BWP7T $T=704360 429400 1 0 $X=704070 $Y=425190
X1266 118 546 3 1 556 DFQD0BWP7T $T=704920 390200 1 0 $X=704630 $Y=385990
X1267 118 545 3 1 562 DFQD0BWP7T $T=704920 398040 0 0 $X=704630 $Y=397805
X1268 118 541 3 1 538 DFQD0BWP7T $T=716680 452920 1 180 $X=705750 $Y=452685
X1269 118 548 3 1 564 DFQD0BWP7T $T=707160 413720 0 0 $X=706870 $Y=413485
X1270 118 549 3 1 566 DFQD0BWP7T $T=707720 437240 0 0 $X=707430 $Y=437005
X1271 118 547 3 1 555 DFQD0BWP7T $T=727880 374520 1 180 $X=716950 $Y=374285
X1272 118 561 3 1 554 DFQD0BWP7T $T=729000 452920 1 180 $X=718070 $Y=452685
X1273 210 580 3 1 570 DFQD0BWP7T $T=738520 366680 1 180 $X=727590 $Y=366445
X1274 118 589 3 1 557 DFQD0BWP7T $T=738520 382360 1 180 $X=727590 $Y=382125
X1275 118 572 3 1 583 DFQD0BWP7T $T=738520 398040 0 180 $X=727590 $Y=393830
X1276 118 571 3 1 587 DFQD0BWP7T $T=738520 413720 0 180 $X=727590 $Y=409510
X1277 118 590 3 1 581 DFQD0BWP7T $T=738520 421560 1 180 $X=727590 $Y=421325
X1278 118 591 3 1 586 DFQD0BWP7T $T=738520 437240 1 180 $X=727590 $Y=437005
X1279 118 582 3 1 575 DFQD0BWP7T $T=738520 452920 0 180 $X=727590 $Y=448710
X1280 118 584 3 1 576 DFQD0BWP7T $T=738520 468600 0 180 $X=727590 $Y=464390
X1281 118 565 3 1 228 DFQD0BWP7T $T=738520 476440 1 180 $X=727590 $Y=476205
X1282 94 3 1 312 327 331 NR3D0BWP7T $T=511720 421560 1 0 $X=511430 $Y=417350
X1283 430 3 1 130 125 425 NR3D0BWP7T $T=598520 382360 1 0 $X=598230 $Y=378150
X1284 309 1 417 401 312 3 AOI21D2BWP7T $T=587880 437240 0 180 $X=582550 $Y=433030
X1285 73 277 271 275 3 1 AOI21D0BWP7T $T=479800 452920 1 180 $X=476710 $Y=452685
X1286 321 310 93 92 3 1 AOI21D0BWP7T $T=512280 468600 1 180 $X=509190 $Y=468365
X1287 275 319 316 324 3 1 AOI21D0BWP7T $T=510600 460760 1 0 $X=510310 $Y=456550
X1288 303 347 312 94 3 1 AOI21D0BWP7T $T=536360 413720 0 0 $X=536070 $Y=413485
X1289 366 379 394 395 3 1 AOI21D0BWP7T $T=562680 421560 0 0 $X=562390 $Y=421325
X1290 410 407 406 381 3 1 AOI21D0BWP7T $T=580040 398040 0 180 $X=576950 $Y=393830
X1291 369 387 303 416 3 1 AOI21D0BWP7T $T=581720 437240 0 0 $X=581430 $Y=437005
X1292 369 416 85 151 3 1 AOI21D0BWP7T $T=587320 437240 0 0 $X=587030 $Y=437005
X1293 385 3 1 370 BUFFD0BWP7T $T=559880 382360 0 0 $X=559590 $Y=382125
X1294 442 3 1 423 BUFFD0BWP7T $T=606920 421560 1 0 $X=606630 $Y=417350
X1295 452 3 1 454 BUFFD0BWP7T $T=622040 468600 0 0 $X=621750 $Y=468365
X1296 131 128 3 1 284 AN2D1BWP7T $T=560440 437240 0 180 $X=557350 $Y=433030
X1297 142 128 3 1 144 AN2D1BWP7T $T=582280 429400 1 0 $X=581990 $Y=425190
X1298 3 1 ICV_61 $T=450120 437240 0 0 $X=449830 $Y=437005
X1299 3 1 ICV_61 $T=479800 398040 0 0 $X=479510 $Y=397805
X1300 3 1 ICV_61 $T=479800 413720 0 0 $X=479510 $Y=413485
X1301 3 1 ICV_61 $T=479800 452920 0 0 $X=479510 $Y=452685
X1302 3 1 ICV_61 $T=521240 366680 0 0 $X=520950 $Y=366445
X1303 3 1 ICV_61 $T=521240 445080 1 0 $X=520950 $Y=440870
X1304 3 1 ICV_61 $T=534120 382360 0 0 $X=533830 $Y=382125
X1305 3 1 ICV_61 $T=605240 382360 0 0 $X=604950 $Y=382125
X1306 3 1 ICV_61 $T=605800 437240 1 0 $X=605510 $Y=433030
X1307 3 1 ICV_61 $T=647240 366680 1 0 $X=646950 $Y=362470
X1308 3 1 ICV_61 $T=666840 382360 0 0 $X=666550 $Y=382125
X1309 3 1 ICV_61 $T=666840 421560 1 0 $X=666550 $Y=417350
X1310 3 1 ICV_61 $T=678040 374520 1 0 $X=677750 $Y=370310
X1311 3 1 ICV_61 $T=689240 437240 0 0 $X=688950 $Y=437005
X1312 3 1 ICV_61 $T=689800 405880 0 0 $X=689510 $Y=405645
X1313 3 1 ICV_61 $T=702120 358840 0 0 $X=701830 $Y=358605
X1314 147 3 418 440 1 421 410 OAI211D0BWP7T $T=606360 390200 1 180 $X=602710 $Y=389965
X1315 433 3 143 149 1 127 442 OAI211D0BWP7T $T=609160 421560 1 0 $X=608870 $Y=417350
X1316 34 250 3 1 23 DFQD1BWP7T $T=468040 421560 1 180 $X=457110 $Y=421325
X1317 34 270 3 1 58 DFQD1BWP7T $T=477000 445080 0 180 $X=466070 $Y=440870
X1318 34 296 3 1 256 DFQD1BWP7T $T=503320 437240 0 180 $X=492390 $Y=433030
X1319 34 304 3 1 246 DFQD1BWP7T $T=506680 421560 1 180 $X=495750 $Y=421325
X1320 34 359 3 1 354 DFQD1BWP7T $T=541960 429400 1 0 $X=541670 $Y=425190
X1321 34 360 3 1 377 DFQD1BWP7T $T=545320 390200 1 0 $X=545030 $Y=385990
X1322 34 370 3 1 382 DFQD1BWP7T $T=548120 398040 0 0 $X=547830 $Y=397805
X1323 118 439 3 1 446 DFQD1BWP7T $T=601320 413720 1 0 $X=601030 $Y=409510
X1324 118 487 3 1 187 DFQD1BWP7T $T=654520 460760 0 180 $X=643590 $Y=456550
X1325 118 502 3 1 208 DFQD1BWP7T $T=683080 484280 0 180 $X=672150 $Y=480070
X1326 262 255 54 52 46 3 1 XNR4D0BWP7T $T=470280 452920 1 180 $X=457110 $Y=452685
X1327 400 431 432 429 155 3 1 XNR4D0BWP7T $T=589560 452920 0 0 $X=589270 $Y=452685
X1328 432 437 159 444 447 3 1 XNR4D0BWP7T $T=599640 460760 1 0 $X=599350 $Y=456550
X1329 377 130 3 1 BUFFD12BWP7T $T=558200 374520 1 0 $X=557910 $Y=370310
X1330 393 438 160 443 448 3 1 XOR4D0BWP7T $T=599640 476440 1 0 $X=599350 $Y=472230
X1331 120 3 1 112 CKND1BWP7T $T=547000 445080 0 0 $X=546710 $Y=444845
X1332 141 3 1 402 CKND1BWP7T $T=621480 445080 0 180 $X=619510 $Y=440870
X1333 149 3 1 441 CKND1BWP7T $T=622040 390200 1 0 $X=621750 $Y=385990
X1334 149 418 3 1 BUFFD1P5BWP7T $T=618680 390200 0 0 $X=618390 $Y=389965
X1335 450 166 3 1 BUFFD1P5BWP7T $T=621480 468600 1 0 $X=621190 $Y=464390
X1336 445 190 3 1 BUFFD1P5BWP7T $T=643320 390200 0 0 $X=643030 $Y=389965
X1337 394 402 1 383 3 354 307 AOI22D1BWP7T $T=570520 437240 0 180 $X=566310 $Y=433030
X1338 130 3 1 127 INVD3BWP7T $T=570520 382360 1 180 $X=566870 $Y=382125
X1339 62 3 1 51 CKBD1BWP7T $T=468040 484280 0 180 $X=465510 $Y=480070
X1340 347 3 1 95 CKBD1BWP7T $T=537480 405880 1 180 $X=534950 $Y=405645
X1341 386 3 1 134 CKBD1BWP7T $T=560440 358840 0 0 $X=560150 $Y=358605
X1342 461 3 1 175 CKBD1BWP7T $T=632680 468600 0 0 $X=632390 $Y=468365
X1343 453 3 1 178 CKBD1BWP7T $T=636040 468600 1 0 $X=635750 $Y=464390
X1344 464 3 1 470 CKBD1BWP7T $T=636600 460760 1 0 $X=636310 $Y=456550
X1345 462 3 1 181 CKBD1BWP7T $T=639400 358840 0 0 $X=639110 $Y=358605
X1346 459 3 1 171 CKBD1BWP7T $T=641080 390200 0 0 $X=640790 $Y=389965
X1347 467 3 1 202 CKBD1BWP7T $T=651720 390200 0 0 $X=651430 $Y=389965
X1348 201 195 1 3 195 196 194 MAOI22D0BWP7T $T=652280 484280 0 180 $X=648070 $Y=480070
X1349 484 203 1 3 203 495 184 MAOI22D0BWP7T $T=664600 366680 1 180 $X=660390 $Y=366445
X1350 529 203 1 3 203 517 516 MAOI22D0BWP7T $T=694840 366680 0 180 $X=690630 $Y=362470
X1351 555 203 1 3 203 547 220 MAOI22D0BWP7T $T=711080 374520 0 180 $X=706870 $Y=370310
X1352 570 203 1 3 203 580 223 MAOI22D0BWP7T $T=721160 366680 0 0 $X=720870 $Y=366445
X1353 31 20 41 8 33 3 1 OAI31D1BWP7T $T=457960 429400 0 180 $X=453750 $Y=425190
X1354 125 127 350 123 124 3 1 OAI31D1BWP7T $T=554280 374520 1 0 $X=553990 $Y=370310
X1355 130 133 386 123 124 3 1 OAI31D1BWP7T $T=565480 358840 0 0 $X=565190 $Y=358605
X1356 112 396 400 297 404 3 1 OAI31D1BWP7T $T=566600 445080 0 0 $X=566310 $Y=444845
X1357 418 143 372 147 124 3 1 OAI31D1BWP7T $T=596280 374520 0 180 $X=592070 $Y=370310
X1358 113 449 437 332 451 3 1 OAI31D1BWP7T $T=620920 452920 1 0 $X=620630 $Y=448710
X1359 141 125 455 127 124 3 1 OAI31D1BWP7T $T=626520 429400 1 180 $X=622310 $Y=429165
X1360 430 441 459 421 124 3 1 OAI31D1BWP7T $T=628200 390200 1 0 $X=627910 $Y=385990
X1361 149 147 173 421 124 3 1 OAI31D1BWP7T $T=630440 366680 1 0 $X=630150 $Y=362470
X1362 149 147 462 421 124 3 1 OAI31D1BWP7T $T=636040 374520 0 180 $X=631830 $Y=370310
X1363 309 310 273 1 3 275 OA21D0BWP7T $T=505560 460760 1 180 $X=501910 $Y=460525
X1364 415 417 434 1 3 439 OA21D0BWP7T $T=599080 405880 0 0 $X=598790 $Y=405645
X1365 12 19 24 29 39 1 3 AOI22D0BWP7T $T=451240 413720 1 0 $X=450950 $Y=409510
X1366 45 248 44 28 38 1 3 AOI22D0BWP7T $T=458520 366680 0 180 $X=454870 $Y=362470
X1367 263 253 23 44 39 1 3 AOI22D0BWP7T $T=471400 429400 0 180 $X=467750 $Y=425190
X1368 45 264 44 265 269 1 3 AOI22D0BWP7T $T=469720 366680 0 0 $X=469430 $Y=366445
X1369 6 261 44 257 265 1 3 AOI22D0BWP7T $T=470280 382360 1 0 $X=469990 $Y=378150
X1370 26 259 44 268 257 1 3 AOI22D0BWP7T $T=470280 390200 1 0 $X=469990 $Y=385990
X1371 53 258 44 263 268 1 3 AOI22D0BWP7T $T=470280 405880 1 0 $X=469990 $Y=401670
X1372 72 280 44 269 74 1 3 AOI22D0BWP7T $T=479800 358840 0 0 $X=479510 $Y=358605
X1373 282 274 11 29 39 1 3 AOI22D0BWP7T $T=483160 413720 0 180 $X=479510 $Y=409510
X1374 26 281 44 272 288 1 3 AOI22D0BWP7T $T=480360 390200 1 0 $X=480070 $Y=385990
X1375 53 276 44 282 272 1 3 AOI22D0BWP7T $T=482600 405880 1 0 $X=482310 $Y=401670
X1376 290 289 256 44 39 1 3 AOI22D0BWP7T $T=486520 413720 0 180 $X=482870 $Y=409510
X1377 315 298 246 44 39 1 3 AOI22D0BWP7T $T=498840 421560 0 180 $X=495190 $Y=417350
X1378 6 300 44 288 90 1 3 AOI22D0BWP7T $T=498840 374520 1 0 $X=498550 $Y=370310
X1379 53 301 44 290 328 1 3 AOI22D0BWP7T $T=503320 398040 0 0 $X=503030 $Y=397805
X1380 6 317 44 323 325 1 3 AOI22D0BWP7T $T=510600 374520 1 0 $X=510310 $Y=370310
X1381 53 320 44 315 329 1 3 AOI22D0BWP7T $T=512280 405880 0 0 $X=511990 $Y=405645
X1382 26 308 44 328 323 1 3 AOI22D0BWP7T $T=517880 390200 1 180 $X=514230 $Y=389965
X1383 6 334 44 333 101 1 3 AOI22D0BWP7T $T=525160 382360 0 180 $X=521510 $Y=378150
X1384 26 336 44 329 333 1 3 AOI22D0BWP7T $T=525160 390200 1 180 $X=521510 $Y=389965
X1385 45 337 44 325 109 1 3 AOI22D0BWP7T $T=528520 366680 0 180 $X=524870 $Y=362470
X1386 479 474 187 151 182 1 3 AOI22D0BWP7T $T=646120 445080 1 180 $X=642470 $Y=444845
X1387 193 477 151 476 475 1 3 AOI22D0BWP7T $T=648360 382360 0 180 $X=644710 $Y=378150
X1388 191 478 151 475 484 1 3 AOI22D0BWP7T $T=646680 366680 0 0 $X=646390 $Y=366445
X1389 482 485 151 479 481 1 3 AOI22D0BWP7T $T=651160 429400 1 180 $X=647510 $Y=429165
X1390 491 486 197 151 182 1 3 AOI22D0BWP7T $T=652280 452920 0 180 $X=648630 $Y=448710
X1391 483 493 151 488 476 1 3 AOI22D0BWP7T $T=654520 405880 0 180 $X=650870 $Y=401670
X1392 480 494 151 481 488 1 3 AOI22D0BWP7T $T=654520 413720 1 180 $X=650870 $Y=413485
X1393 482 496 151 491 509 1 3 AOI22D0BWP7T $T=660680 437240 0 0 $X=660390 $Y=437005
X1394 513 498 204 151 182 1 3 AOI22D0BWP7T $T=664040 460760 1 180 $X=660390 $Y=460525
X1395 512 510 209 151 182 1 3 AOI22D0BWP7T $T=676360 468600 0 180 $X=672710 $Y=464390
X1396 480 507 151 509 514 1 3 AOI22D0BWP7T $T=673560 413720 0 0 $X=673270 $Y=413485
X1397 482 508 151 513 515 1 3 AOI22D0BWP7T $T=674120 445080 1 0 $X=673830 $Y=440870
X1398 483 511 151 514 214 1 3 AOI22D0BWP7T $T=680840 398040 1 0 $X=680550 $Y=393830
X1399 193 506 151 520 526 1 3 AOI22D0BWP7T $T=681960 390200 1 0 $X=681670 $Y=385990
X1400 480 527 151 515 525 1 3 AOI22D0BWP7T $T=687000 421560 1 0 $X=686710 $Y=417350
X1401 482 531 151 512 533 1 3 AOI22D0BWP7T $T=688120 445080 0 0 $X=687830 $Y=444845
X1402 191 522 151 526 529 1 3 AOI22D0BWP7T $T=692600 374520 0 180 $X=688950 $Y=370310
X1403 480 528 151 533 534 1 3 AOI22D0BWP7T $T=691480 437240 1 0 $X=691190 $Y=433030
X1404 483 542 151 525 218 1 3 AOI22D0BWP7T $T=706040 382360 0 180 $X=702390 $Y=378150
X1405 483 532 151 534 520 1 3 AOI22D0BWP7T $T=702680 413720 1 0 $X=702390 $Y=409510
X1406 482 539 151 538 543 1 3 AOI22D0BWP7T $T=702680 437240 0 0 $X=702390 $Y=437005
X1407 538 537 215 151 182 1 3 AOI22D0BWP7T $T=702680 460760 0 0 $X=702390 $Y=460525
X1408 554 552 219 151 182 1 3 AOI22D0BWP7T $T=711640 468600 0 180 $X=707990 $Y=464390
X1409 483 550 151 556 226 1 3 AOI22D0BWP7T $T=709400 382360 0 0 $X=709110 $Y=382125
X1410 480 553 151 543 556 1 3 AOI22D0BWP7T $T=710520 413720 1 0 $X=710230 $Y=409510
X1411 191 559 151 557 555 1 3 AOI22D0BWP7T $T=715000 374520 1 180 $X=711350 $Y=374285
X1412 482 558 151 554 566 1 3 AOI22D0BWP7T $T=712760 452920 1 0 $X=712470 $Y=448710
X1413 480 560 151 566 587 1 3 AOI22D0BWP7T $T=716680 429400 1 0 $X=716390 $Y=425190
X1414 191 563 151 573 570 1 3 AOI22D0BWP7T $T=719480 358840 0 0 $X=719190 $Y=358605
X1415 482 568 151 228 575 1 3 AOI22D0BWP7T $T=720040 460760 0 0 $X=719750 $Y=460525
X1416 576 229 227 151 182 1 3 AOI22D0BWP7T $T=723400 476440 1 180 $X=719750 $Y=476205
X1417 193 569 151 583 573 1 3 AOI22D0BWP7T $T=721720 382360 0 0 $X=721430 $Y=382125
X1418 483 578 151 581 562 1 3 AOI22D0BWP7T $T=722840 421560 1 0 $X=722550 $Y=417350
X1419 480 579 151 575 564 1 3 AOI22D0BWP7T $T=726200 437240 0 180 $X=722550 $Y=433030
X1420 193 567 151 562 557 1 3 AOI22D0BWP7T $T=723960 398040 1 0 $X=723670 $Y=393830
X1421 483 574 151 564 230 1 3 AOI22D0BWP7T $T=723960 405880 0 0 $X=723670 $Y=405645
X1422 480 585 151 586 581 1 3 AOI22D0BWP7T $T=726200 429400 0 0 $X=725910 $Y=429165
X1423 483 577 151 587 583 1 3 AOI22D0BWP7T $T=735160 405880 1 0 $X=734870 $Y=401670
X1424 482 588 151 576 586 1 3 AOI22D0BWP7T $T=738520 460760 0 180 $X=734870 $Y=456550
X1425 3 1 ICV_41 $T=450120 398040 1 0 $X=449830 $Y=393830
X1426 3 1 ICV_41 $T=475880 476440 0 0 $X=475590 $Y=476205
X1427 3 1 ICV_41 $T=476440 366680 1 0 $X=476150 $Y=362470
X1428 3 1 ICV_41 $T=477000 445080 1 0 $X=476710 $Y=440870
X1429 3 1 ICV_41 $T=517880 421560 0 0 $X=517590 $Y=421325
X1430 3 1 ICV_41 $T=517880 468600 1 0 $X=517590 $Y=464390
X1431 3 1 ICV_41 $T=518440 476440 0 0 $X=518150 $Y=476205
X1432 3 1 ICV_41 $T=519000 460760 1 0 $X=518710 $Y=456550
X1433 3 1 ICV_41 $T=559880 484280 1 0 $X=559590 $Y=480070
X1434 3 1 ICV_41 $T=560440 476440 0 0 $X=560150 $Y=476205
X1435 3 1 ICV_41 $T=576120 452920 0 0 $X=575830 $Y=452685
X1436 3 1 ICV_41 $T=602440 437240 0 0 $X=602150 $Y=437005
X1437 3 1 ICV_41 $T=602440 452920 0 0 $X=602150 $Y=452685
X1438 3 1 ICV_41 $T=618120 460760 1 0 $X=617830 $Y=456550
X1439 3 1 ICV_41 $T=660120 429400 1 0 $X=659830 $Y=425190
X1440 3 1 ICV_41 $T=671880 476440 1 0 $X=671590 $Y=472230
X1441 3 1 ICV_41 $T=702120 468600 0 0 $X=701830 $Y=468365
X1442 3 1 ICV_41 $T=720040 460760 1 0 $X=719750 $Y=456550
X1443 3 1 ICV_41 $T=729000 374520 1 0 $X=728710 $Y=370310
X1444 3 1 ICV_41 $T=729000 452920 0 0 $X=728710 $Y=452685
X1445 3 1 ICV_37 $T=450120 374520 0 0 $X=449830 $Y=374285
X1446 3 1 ICV_37 $T=450120 390200 1 0 $X=449830 $Y=385990
X1447 3 1 ICV_37 $T=450120 429400 1 0 $X=449830 $Y=425190
X1448 3 1 ICV_37 $T=480920 468600 1 0 $X=480630 $Y=464390
X1449 3 1 ICV_37 $T=487640 405880 0 0 $X=487350 $Y=405645
X1450 3 1 ICV_37 $T=517880 382360 1 0 $X=517590 $Y=378150
X1451 3 1 ICV_37 $T=519000 484280 1 0 $X=518710 $Y=480070
X1452 3 1 ICV_37 $T=529640 413720 0 0 $X=529350 $Y=413485
X1453 3 1 ICV_37 $T=546440 374520 1 0 $X=546150 $Y=370310
X1454 3 1 ICV_37 $T=552040 398040 1 0 $X=551750 $Y=393830
X1455 3 1 ICV_37 $T=576120 390200 1 0 $X=575830 $Y=385990
X1456 3 1 ICV_37 $T=576120 421560 1 0 $X=575830 $Y=417350
X1457 3 1 ICV_37 $T=618120 374520 0 0 $X=617830 $Y=374285
X1458 3 1 ICV_37 $T=618120 382360 1 0 $X=617830 $Y=378150
X1459 3 1 ICV_37 $T=618120 437240 0 0 $X=617830 $Y=437005
X1460 3 1 ICV_37 $T=618120 452920 0 0 $X=617830 $Y=452685
X1461 3 1 ICV_37 $T=618120 468600 1 0 $X=617830 $Y=464390
X1462 3 1 ICV_37 $T=626520 429400 0 0 $X=626230 $Y=429165
X1463 3 1 ICV_37 $T=636040 358840 0 0 $X=635750 $Y=358605
X1464 3 1 ICV_37 $T=637720 390200 0 0 $X=637430 $Y=389965
X1465 3 1 ICV_37 $T=637720 452920 0 0 $X=637430 $Y=452685
X1466 3 1 ICV_37 $T=655640 413720 1 0 $X=655350 $Y=409510
X1467 3 1 ICV_37 $T=660120 382360 0 0 $X=659830 $Y=382125
X1468 3 1 ICV_37 $T=660120 413720 1 0 $X=659830 $Y=409510
X1469 3 1 ICV_37 $T=660120 421560 1 0 $X=659830 $Y=417350
X1470 3 1 ICV_37 $T=677480 460760 0 0 $X=677190 $Y=460525
X1471 3 1 ICV_37 $T=688120 437240 1 0 $X=687830 $Y=433030
X1472 3 1 ICV_37 $T=716120 358840 0 0 $X=715830 $Y=358605
X1473 3 1 ICV_37 $T=720040 405880 0 0 $X=719750 $Y=405645
X1474 3 1 ICV_37 $T=720040 445080 0 0 $X=719750 $Y=444845
X1475 3 1 ICV_37 $T=731800 405880 1 0 $X=731510 $Y=401670
X1476 3 1 ICV_60 $T=450120 366680 1 0 $X=449830 $Y=362470
X1477 3 1 ICV_60 $T=454600 413720 1 0 $X=454310 $Y=409510
X1478 3 1 ICV_60 $T=468040 460760 0 0 $X=467750 $Y=460525
X1479 3 1 ICV_60 $T=470280 452920 0 0 $X=469990 $Y=452685
X1480 3 1 ICV_60 $T=470840 437240 1 0 $X=470550 $Y=433030
X1481 3 1 ICV_60 $T=477000 484280 1 0 $X=476710 $Y=480070
X1482 3 1 ICV_60 $T=492120 398040 0 0 $X=491830 $Y=397805
X1483 3 1 ICV_60 $T=496600 452920 0 0 $X=496310 $Y=452685
X1484 3 1 ICV_60 $T=501080 382360 1 0 $X=500790 $Y=378150
X1485 3 1 ICV_60 $T=515640 405880 0 0 $X=515350 $Y=405645
X1486 3 1 ICV_60 $T=536920 468600 0 0 $X=536630 $Y=468365
X1487 3 1 ICV_60 $T=548680 452920 1 0 $X=548390 $Y=448710
X1488 3 1 ICV_60 $T=585080 468600 1 0 $X=584790 $Y=464390
X1489 3 1 ICV_60 $T=585080 484280 1 0 $X=584790 $Y=480070
X1490 3 1 ICV_60 $T=627080 374520 1 0 $X=626790 $Y=370310
X1491 3 1 ICV_60 $T=702120 374520 1 0 $X=701830 $Y=370310
X1492 3 1 ICV_60 $T=702120 405880 1 0 $X=701830 $Y=401670
X1493 3 1 ICV_60 $T=702120 413720 0 0 $X=701830 $Y=413485
X1494 3 1 ICV_60 $T=715000 460760 0 0 $X=714710 $Y=460525
X1495 3 1 ICV_43 $T=450120 445080 1 0 $X=449830 $Y=440870
X1496 3 1 ICV_43 $T=534120 382360 1 0 $X=533830 $Y=378150
X1497 3 1 ICV_43 $T=534120 413720 1 0 $X=533830 $Y=409510
X1498 3 1 ICV_43 $T=545320 413720 1 0 $X=545030 $Y=409510
X1499 3 1 ICV_43 $T=554840 437240 1 0 $X=554550 $Y=433030
X1500 3 1 ICV_43 $T=561000 366680 0 0 $X=560710 $Y=366445
X1501 3 1 ICV_43 $T=561560 437240 0 0 $X=561270 $Y=437005
X1502 3 1 ICV_43 $T=576120 452920 1 0 $X=575830 $Y=448710
X1503 3 1 ICV_43 $T=581720 405880 0 0 $X=581430 $Y=405645
X1504 3 1 ICV_43 $T=584520 437240 0 0 $X=584230 $Y=437005
X1505 3 1 ICV_43 $T=624280 468600 0 0 $X=623990 $Y=468365
X1506 3 1 ICV_43 $T=627080 405880 1 0 $X=626790 $Y=401670
X1507 3 1 ICV_43 $T=633240 468600 1 0 $X=632950 $Y=464390
X1508 3 1 ICV_43 $T=685880 429400 1 0 $X=685590 $Y=425190
X1509 3 1 ICV_43 $T=702120 390200 1 0 $X=701830 $Y=385990
X1510 3 1 ICV_43 $T=702120 398040 0 0 $X=701830 $Y=397805
X1511 3 1 ICV_43 $T=720040 421560 1 0 $X=719750 $Y=417350
X1512 3 1 ICV_43 $T=720040 437240 1 0 $X=719750 $Y=433030
X1513 3 1 ICV_43 $T=725080 452920 1 0 $X=724790 $Y=448710
X1514 3 1 ICV_52 $T=470280 413720 1 0 $X=469990 $Y=409510
X1515 3 1 ICV_52 $T=492120 366680 1 0 $X=491830 $Y=362470
X1516 3 1 ICV_52 $T=492120 421560 0 0 $X=491830 $Y=421325
X1517 3 1 ICV_52 $T=505000 398040 1 0 $X=504710 $Y=393830
X1518 3 1 ICV_52 $T=517880 390200 0 0 $X=517590 $Y=389965
X1519 3 1 ICV_52 $T=529080 382360 0 0 $X=528790 $Y=382125
X1520 3 1 ICV_52 $T=529080 484280 1 0 $X=528790 $Y=480070
X1521 3 1 ICV_52 $T=562680 437240 1 0 $X=562390 $Y=433030
X1522 3 1 ICV_52 $T=564360 452920 1 0 $X=564070 $Y=448710
X1523 3 1 ICV_52 $T=571080 468600 0 0 $X=570790 $Y=468365
X1524 3 1 ICV_52 $T=576120 358840 0 0 $X=575830 $Y=358605
X1525 3 1 ICV_52 $T=603000 445080 1 0 $X=602710 $Y=440870
X1526 3 1 ICV_52 $T=613080 398040 0 0 $X=612790 $Y=397805
X1527 3 1 ICV_52 $T=613080 452920 1 0 $X=612790 $Y=448710
X1528 3 1 ICV_52 $T=618120 429400 1 0 $X=617830 $Y=425190
X1529 3 1 ICV_52 $T=618120 468600 0 0 $X=617830 $Y=468365
X1530 3 1 ICV_52 $T=626520 366680 1 0 $X=626230 $Y=362470
X1531 3 1 ICV_52 $T=641080 382360 1 0 $X=640790 $Y=378150
X1532 3 1 ICV_52 $T=655080 445080 0 0 $X=654790 $Y=444845
X1533 3 1 ICV_52 $T=669080 405880 1 0 $X=668790 $Y=401670
X1534 3 1 ICV_52 $T=678040 452920 1 0 $X=677750 $Y=448710
X1535 3 1 ICV_52 $T=697080 374520 1 0 $X=696790 $Y=370310
X1536 3 1 ICV_52 $T=702120 452920 0 0 $X=701830 $Y=452685
X1537 8 1 27 40 3 NR2XD0BWP7T $T=452920 476440 0 0 $X=452630 $Y=476205
X1538 3 1 ICV_38 $T=486520 358840 0 0 $X=486230 $Y=358605
X1539 3 1 ICV_38 $T=486520 366680 0 0 $X=486230 $Y=366445
X1540 3 1 ICV_38 $T=486520 382360 1 0 $X=486230 $Y=378150
X1541 3 1 ICV_38 $T=486520 413720 1 0 $X=486230 $Y=409510
X1542 3 1 ICV_38 $T=486520 429400 1 0 $X=486230 $Y=425190
X1543 3 1 ICV_38 $T=486520 437240 1 0 $X=486230 $Y=433030
X1544 3 1 ICV_38 $T=486520 445080 0 0 $X=486230 $Y=444845
X1545 3 1 ICV_38 $T=486520 468600 1 0 $X=486230 $Y=464390
X1546 3 1 ICV_38 $T=486520 476440 1 0 $X=486230 $Y=472230
X1547 3 1 ICV_38 $T=528520 382360 1 0 $X=528230 $Y=378150
X1548 3 1 ICV_38 $T=528520 437240 1 0 $X=528230 $Y=433030
X1549 3 1 ICV_38 $T=528520 460760 0 0 $X=528230 $Y=460525
X1550 3 1 ICV_38 $T=570520 366680 0 0 $X=570230 $Y=366445
X1551 3 1 ICV_38 $T=570520 374520 1 0 $X=570230 $Y=370310
X1552 3 1 ICV_38 $T=570520 382360 0 0 $X=570230 $Y=382125
X1553 3 1 ICV_38 $T=570520 421560 0 0 $X=570230 $Y=421325
X1554 3 1 ICV_38 $T=570520 429400 1 0 $X=570230 $Y=425190
X1555 3 1 ICV_38 $T=570520 437240 1 0 $X=570230 $Y=433030
X1556 3 1 ICV_38 $T=570520 445080 0 0 $X=570230 $Y=444845
X1557 3 1 ICV_38 $T=570520 452920 1 0 $X=570230 $Y=448710
X1558 3 1 ICV_38 $T=570520 460760 1 0 $X=570230 $Y=456550
X1559 3 1 ICV_38 $T=570520 476440 1 0 $X=570230 $Y=472230
X1560 3 1 ICV_38 $T=612520 358840 0 0 $X=612230 $Y=358605
X1561 3 1 ICV_38 $T=612520 374520 0 0 $X=612230 $Y=374285
X1562 3 1 ICV_38 $T=612520 382360 1 0 $X=612230 $Y=378150
X1563 3 1 ICV_38 $T=612520 460760 1 0 $X=612230 $Y=456550
X1564 3 1 ICV_38 $T=612520 476440 1 0 $X=612230 $Y=472230
X1565 3 1 ICV_38 $T=654520 382360 1 0 $X=654230 $Y=378150
X1566 3 1 ICV_38 $T=654520 460760 1 0 $X=654230 $Y=456550
X1567 3 1 ICV_38 $T=696520 358840 0 0 $X=696230 $Y=358605
X1568 3 1 ICV_38 $T=696520 374520 0 0 $X=696230 $Y=374285
X1569 3 1 ICV_38 $T=696520 382360 0 0 $X=696230 $Y=382125
X1570 3 1 ICV_38 $T=696520 398040 0 0 $X=696230 $Y=397805
X1571 3 1 ICV_38 $T=696520 445080 0 0 $X=696230 $Y=444845
X1572 3 1 ICV_38 $T=696520 460760 1 0 $X=696230 $Y=456550
X1573 3 1 ICV_38 $T=696520 476440 1 0 $X=696230 $Y=472230
X1574 3 1 ICV_45 $T=463560 437240 0 0 $X=463270 $Y=437005
X1575 3 1 ICV_45 $T=492120 484280 1 0 $X=491830 $Y=480070
X1576 3 1 ICV_45 $T=502760 413720 0 0 $X=502470 $Y=413485
X1577 3 1 ICV_45 $T=534120 366680 0 0 $X=533830 $Y=366445
X1578 3 1 ICV_45 $T=534120 460760 1 0 $X=533830 $Y=456550
X1579 3 1 ICV_45 $T=544200 468600 0 0 $X=543910 $Y=468365
X1580 3 1 ICV_45 $T=547000 452920 0 0 $X=546710 $Y=452685
X1581 3 1 ICV_45 $T=548120 366680 1 0 $X=547830 $Y=362470
X1582 3 1 ICV_45 $T=576120 405880 1 0 $X=575830 $Y=401670
X1583 3 1 ICV_45 $T=576120 445080 1 0 $X=575830 $Y=440870
X1584 3 1 ICV_45 $T=585640 374520 0 0 $X=585350 $Y=374285
X1585 3 1 ICV_45 $T=586200 452920 1 0 $X=585910 $Y=448710
X1586 3 1 ICV_45 $T=588440 421560 0 0 $X=588150 $Y=421325
X1587 3 1 ICV_45 $T=589560 366680 0 0 $X=589270 $Y=366445
X1588 3 1 ICV_45 $T=590120 460760 0 0 $X=589830 $Y=460525
X1589 3 1 ICV_45 $T=624840 437240 1 0 $X=624550 $Y=433030
X1590 3 1 ICV_45 $T=624840 460760 0 0 $X=624550 $Y=460525
X1591 3 1 ICV_45 $T=628760 413720 1 0 $X=628470 $Y=409510
X1592 3 1 ICV_45 $T=714440 476440 1 0 $X=714150 $Y=472230
X1593 3 1 ICV_45 $T=715000 445080 1 0 $X=714710 $Y=440870
X1594 354 312 3 1 INVD2P5BWP7T $T=545320 421560 0 180 $X=542230 $Y=417350
X1595 430 147 3 1 INVD2P5BWP7T $T=611960 374520 0 180 $X=608870 $Y=370310
X1596 465 97 3 1 INVD2P5BWP7T $T=638280 382360 1 0 $X=637990 $Y=378150
X1597 446 3 1 143 BUFFD3BWP7T $T=610280 429400 1 180 $X=606070 $Y=429165
X1598 350 3 1 311 BUFFD1BWP7T $T=539160 382360 0 180 $X=536630 $Y=378150
X1599 372 3 1 121 BUFFD1BWP7T $T=552600 374520 0 180 $X=550070 $Y=370310
X1600 455 3 1 466 BUFFD1BWP7T $T=634360 460760 1 0 $X=634070 $Y=456550
X1601 143 150 3 1 156 467 IAO21D0BWP7T $T=634360 390200 0 0 $X=634070 $Y=389965
X1602 369 344 303 1 3 345 AN3D1BWP7T $T=559880 445080 1 180 $X=556230 $Y=444845
X1603 216 1 118 3 CKND12BWP7T $T=692040 484280 0 180 $X=682790 $Y=480070
X1604 118 424 149 3 1 DFQD2BWP7T $T=589000 413720 0 0 $X=588710 $Y=413485
X1605 118 426 430 3 1 DFQD2BWP7T $T=600200 398040 1 0 $X=599910 $Y=393830
X1606 118 490 197 3 1 DFQD2BWP7T $T=671880 476440 0 180 $X=660390 $Y=472230
X1607 118 536 215 3 1 DFQD2BWP7T $T=696520 476440 0 180 $X=685030 $Y=472230
X1608 118 551 219 3 1 DFQD2BWP7T $T=713880 476440 1 180 $X=702390 $Y=476205
X1609 29 3 1 151 BUFFD5BWP7T $T=588440 398040 1 0 $X=588150 $Y=393830
X1610 171 170 166 3 1 ND2D2BWP7T $T=631000 468600 1 180 $X=626790 $Y=468365
X1611 460 177 166 3 1 ND2D2BWP7T $T=639960 476440 1 180 $X=635750 $Y=476205
X1612 169 183 466 3 1 ND2D2BWP7T $T=638840 484280 1 0 $X=638550 $Y=480070
X1613 456 188 473 3 1 ND2D2BWP7T $T=642200 413720 0 0 $X=641910 $Y=413485
X1614 460 192 470 3 1 ND2D2BWP7T $T=645000 468600 0 0 $X=644710 $Y=468365
X1615 107 199 470 3 1 ND2D2BWP7T $T=648360 476440 1 0 $X=648070 $Y=472230
X1616 91 39 311 3 1 ND2D1P5BWP7T $T=501640 366680 0 0 $X=501350 $Y=366445
X1617 97 53 311 3 1 ND2D1P5BWP7T $T=516200 382360 0 0 $X=515910 $Y=382125
X1618 107 6 311 3 1 ND2D1P5BWP7T $T=525160 374520 0 180 $X=520950 $Y=370310
X1619 122 26 311 3 1 ND2D1P5BWP7T $T=551480 374520 1 180 $X=547270 $Y=374285
X1620 441 150 147 3 1 ND2D1P5BWP7T $T=621480 374520 0 0 $X=621190 $Y=374285
X1621 97 176 454 3 1 ND2D1P5BWP7T $T=638840 476440 0 180 $X=634630 $Y=472230
X1622 169 191 190 3 1 ND2D1P5BWP7T $T=643320 366680 1 0 $X=643030 $Y=362470
X1623 181 182 190 3 1 ND2D1P5BWP7T $T=645000 437240 0 0 $X=644710 $Y=437005
X1624 458 480 190 3 1 ND2D1P5BWP7T $T=646120 413720 0 0 $X=645830 $Y=413485
X1625 171 482 190 3 1 ND2D1P5BWP7T $T=646120 445080 1 0 $X=645830 $Y=440870
X1626 107 483 190 3 1 ND2D1P5BWP7T $T=646680 390200 0 0 $X=646390 $Y=389965
X1628 307 3 305 89 1 292 87 OAI211D1BWP7T $T=503320 445080 0 180 $X=499670 $Y=440870
X1629 389 3 352 141 1 ND2D4BWP7T $T=591240 437240 0 0 $X=590950 $Y=437005
X1630 309 1 345 348 3 349 351 AOI211D1BWP7T $T=535240 445080 0 0 $X=534950 $Y=444845
X1631 309 1 383 368 3 355 358 AOI211D1BWP7T $T=561560 437240 1 180 $X=557910 $Y=437005
X1632 381 1 395 413 3 415 143 AOI211D1BWP7T $T=580040 421560 1 0 $X=579750 $Y=417350
X1633 71 27 3 1 BUFFD8BWP7T $T=477560 429400 1 0 $X=477270 $Y=425190
X1634 341 71 3 1 BUFFD8BWP7T $T=528520 437240 0 180 $X=519270 $Y=433030
X1635 65 3 57 63 1 61 ND3D1BWP7T $T=470280 468600 0 180 $X=466630 $Y=464390
X1636 352 3 413 421 1 409 ND3D1BWP7T $T=584520 405880 0 0 $X=584230 $Y=405645
X1637 354 379 1 95 376 3 OAI21D1BWP7T $T=553720 421560 1 0 $X=553430 $Y=417350
X1638 150 421 1 124 165 3 OAI21D1BWP7T $T=622040 366680 0 180 $X=618390 $Y=362470
X1639 139 141 1 124 450 3 OAI21D1BWP7T $T=624840 437240 1 180 $X=621190 $Y=437005
X1640 150 421 1 124 458 3 OAI21D1BWP7T $T=628760 413720 0 180 $X=625110 $Y=409510
X1692 114 119 117 3 1 INR2XD2BWP7T $T=541960 366680 1 0 $X=541670 $Y=362470
X1693 473 180 195 3 1 INR2XD2BWP7T $T=645000 405880 1 0 $X=644710 $Y=401670
X1694 190 202 203 3 1 INR2XD2BWP7T $T=648360 382360 1 0 $X=648070 $Y=378150
X1695 29 44 3 1 BUFFD4BWP7T $T=525720 405880 1 180 $X=520390 $Y=405645
X1696 457 169 3 1 BUFFD4BWP7T $T=629320 366680 1 180 $X=623990 $Y=366445
X1697 3 1 ICV_51 $T=489320 452920 1 0 $X=489030 $Y=448710
X1698 3 1 ICV_51 $T=489320 476440 0 0 $X=489030 $Y=476205
X1699 3 1 ICV_51 $T=531320 421560 0 0 $X=531030 $Y=421325
X1700 3 1 ICV_51 $T=531320 468600 1 0 $X=531030 $Y=464390
X1701 3 1 ICV_51 $T=531320 468600 0 0 $X=531030 $Y=468365
X1702 3 1 ICV_51 $T=531320 476440 1 0 $X=531030 $Y=472230
X1703 3 1 ICV_51 $T=573320 413720 1 0 $X=573030 $Y=409510
X1704 3 1 ICV_51 $T=573320 437240 0 0 $X=573030 $Y=437005
X1705 3 1 ICV_51 $T=573320 484280 1 0 $X=573030 $Y=480070
X1706 3 1 ICV_51 $T=615320 390200 0 0 $X=615030 $Y=389965
X1707 3 1 ICV_51 $T=615320 405880 1 0 $X=615030 $Y=401670
X1708 3 1 ICV_51 $T=615320 421560 0 0 $X=615030 $Y=421325
X1709 3 1 ICV_51 $T=615320 429400 1 0 $X=615030 $Y=425190
X1710 3 1 ICV_51 $T=657320 358840 0 0 $X=657030 $Y=358605
X1711 3 1 ICV_51 $T=657320 366680 0 0 $X=657030 $Y=366445
X1712 3 1 ICV_51 $T=657320 374520 0 0 $X=657030 $Y=374285
X1713 3 1 ICV_51 $T=699320 366680 1 0 $X=699030 $Y=362470
X1714 3 1 ICV_51 $T=699320 405880 1 0 $X=699030 $Y=401670
X1715 3 1 ICV_51 $T=699320 413720 0 0 $X=699030 $Y=413485
X1716 3 1 ICV_51 $T=699320 421560 1 0 $X=699030 $Y=417350
X1717 3 1 ICV_51 $T=699320 437240 1 0 $X=699030 $Y=433030
X1718 85 3 341 139 409 1 OAI21D2BWP7T $T=581720 405880 1 180 $X=576390 $Y=405645
X1719 124 3 122 150 421 1 OAI21D2BWP7T $T=597960 374520 1 0 $X=597670 $Y=370310
X1720 124 3 460 150 421 1 OAI21D2BWP7T $T=627080 398040 1 0 $X=626790 $Y=393830
X1721 141 1 139 94 3 179 NR3D3BWP7T $T=628200 445080 1 0 $X=627910 $Y=440870
X1722 143 150 156 157 1 3 IAO21D2BWP7T $T=603000 374520 1 0 $X=602710 $Y=370310
X1723 149 143 147 124 3 1 145 OA31D0BWP7T $T=589560 366680 1 180 $X=584790 $Y=366445
X1724 430 441 421 124 3 1 465 OA31D0BWP7T $T=631560 382360 1 0 $X=631270 $Y=378150
X1760 3 1 ICV_39 $T=486520 398040 1 0 $X=486230 $Y=393830
X1761 3 1 ICV_39 $T=570520 398040 1 0 $X=570230 $Y=393830
X1762 3 1 ICV_39 $T=570520 460760 0 0 $X=570230 $Y=460525
X1763 3 1 ICV_39 $T=738520 366680 0 0 $X=738230 $Y=366445
X1764 3 1 ICV_39 $T=738520 374520 0 0 $X=738230 $Y=374285
X1765 3 1 ICV_39 $T=738520 382360 0 0 $X=738230 $Y=382125
X1766 3 1 ICV_39 $T=738520 398040 1 0 $X=738230 $Y=393830
X1767 3 1 ICV_39 $T=738520 405880 1 0 $X=738230 $Y=401670
X1768 3 1 ICV_39 $T=738520 413720 1 0 $X=738230 $Y=409510
X1769 3 1 ICV_39 $T=738520 421560 0 0 $X=738230 $Y=421325
X1770 3 1 ICV_39 $T=738520 429400 0 0 $X=738230 $Y=429165
X1771 3 1 ICV_39 $T=738520 437240 1 0 $X=738230 $Y=433030
X1772 3 1 ICV_39 $T=738520 437240 0 0 $X=738230 $Y=437005
X1773 3 1 ICV_39 $T=738520 452920 1 0 $X=738230 $Y=448710
X1774 3 1 ICV_39 $T=738520 460760 1 0 $X=738230 $Y=456550
X1775 3 1 ICV_39 $T=738520 468600 1 0 $X=738230 $Y=464390
X1776 3 1 ICV_39 $T=738520 476440 0 0 $X=738230 $Y=476205
X1777 3 1 ICV_42 $T=492120 476440 0 0 $X=491830 $Y=476205
X1778 3 1 ICV_42 $T=515640 468600 0 0 $X=515350 $Y=468365
X1779 3 1 ICV_42 $T=516200 374520 0 0 $X=515910 $Y=374285
X1780 3 1 ICV_42 $T=587320 445080 0 0 $X=587030 $Y=444845
X1781 3 1 ICV_42 $T=599640 429400 1 0 $X=599350 $Y=425190
X1782 3 1 ICV_42 $T=600200 413720 0 0 $X=599910 $Y=413485
X1783 3 1 ICV_42 $T=618120 476440 1 0 $X=617830 $Y=472230
X1784 3 1 ICV_42 $T=625400 374520 0 0 $X=625110 $Y=374285
X1785 3 1 ICV_42 $T=660120 358840 0 0 $X=659830 $Y=358605
X1786 3 1 ICV_42 $T=660120 374520 0 0 $X=659830 $Y=374285
X1787 3 1 ICV_42 $T=666840 413720 1 0 $X=666550 $Y=409510
X1788 3 1 ICV_42 $T=684200 398040 1 0 $X=683910 $Y=393830
X1789 3 1 ICV_42 $T=684760 366680 0 0 $X=684470 $Y=366445
X1790 3 1 ICV_42 $T=685320 390200 1 0 $X=685030 $Y=385990
X1791 3 1 ICV_42 $T=702120 390200 0 0 $X=701830 $Y=389965
X1792 3 1 ICV_42 $T=726200 445080 0 0 $X=725910 $Y=444845
X1793 3 1 ICV_42 $T=727320 405880 0 0 $X=727030 $Y=405645
X1794 293 65 309 292 312 1 3 314 OA32D0BWP7T $T=501640 452920 0 0 $X=501350 $Y=452685
X1795 130 378 381 127 376 1 3 361 OA32D0BWP7T $T=559880 382360 1 180 $X=553990 $Y=382125
X1796 331 29 3 1 BUFFD6BWP7T $T=520680 421560 1 0 $X=520390 $Y=417350
X1797 371 124 3 1 BUFFD6BWP7T $T=559880 413720 1 0 $X=559590 $Y=409510
X1798 124 3 114 123 125 127 1 OAI31D2BWP7T $T=553160 358840 0 0 $X=552870 $Y=358605
X1799 124 3 136 123 125 127 1 OAI31D2BWP7T $T=570520 366680 1 180 $X=563510 $Y=366445
X1800 124 3 153 147 418 143 1 OAI31D2BWP7T $T=592360 382360 0 0 $X=592070 $Y=382125
X1801 124 3 445 141 130 133 1 OAI31D2BWP7T $T=612520 382360 0 180 $X=605510 $Y=378150
X1802 124 3 453 421 149 147 1 OAI31D2BWP7T $T=625400 421560 0 180 $X=618390 $Y=417350
X1803 124 3 456 147 418 143 1 OAI31D2BWP7T $T=627080 405880 0 180 $X=620070 $Y=401670
X1804 124 3 457 441 430 143 1 OAI31D2BWP7T $T=628200 382360 0 180 $X=621190 $Y=378150
X1805 124 3 461 147 149 143 1 OAI31D2BWP7T $T=634360 421560 0 180 $X=627350 $Y=417350
X1806 124 3 464 141 125 127 1 OAI31D2BWP7T $T=636600 405880 0 180 $X=629590 $Y=401670
X1807 124 3 452 127 141 125 1 OAI31D2BWP7T $T=634920 413720 0 0 $X=634630 $Y=413485
X1808 124 3 473 141 125 127 1 OAI31D2BWP7T $T=643880 405880 0 180 $X=636870 $Y=401670
X1809 130 3 139 125 1 ND2D3BWP7T $T=581720 374520 0 180 $X=576390 $Y=370310
X1810 409 3 107 124 1 ND2D3BWP7T $T=579480 390200 1 0 $X=579190 $Y=385990
X1811 389 3 1 366 CKND0BWP7T $T=578920 437240 1 0 $X=578630 $Y=433030
X1812 418 417 420 309 3 1 424 AO211D0BWP7T $T=584520 421560 0 0 $X=584230 $Y=421325
X1813 125 150 425 423 3 1 397 AO211D0BWP7T $T=590680 382360 1 180 $X=586470 $Y=382125
X1814 430 417 407 309 3 1 426 AO211D0BWP7T $T=592360 405880 1 180 $X=588150 $Y=405645
.ENDS
***************************************
.SUBCKT ICV_56 1 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214
** N=562 EP=212 IP=4154 FDC=10716
*.SEEDPROM
M0 243 41 4 4 N L=1.8e-07 W=5.7e-07 $X=460445 $Y=492465 $D=0
M1 4 41 243 4 N L=1.8e-07 W=5.7e-07 $X=461165 $Y=492465 $D=0
M2 243 41 4 4 N L=1.8e-07 W=5.7e-07 $X=461885 $Y=492465 $D=0
M3 4 41 243 4 N L=1.8e-07 W=5.7e-07 $X=462605 $Y=492465 $D=0
M4 243 41 4 4 N L=1.8e-07 W=5.7e-07 $X=463325 $Y=492465 $D=0
M5 4 41 243 4 N L=1.8e-07 W=5.7e-07 $X=464045 $Y=492465 $D=0
M6 243 41 4 4 N L=1.8e-07 W=5.7e-07 $X=464765 $Y=492465 $D=0
M7 4 37 243 4 N L=1.8e-07 W=5.7e-07 $X=465485 $Y=492465 $D=0
M8 243 37 4 4 N L=1.8e-07 W=5.7e-07 $X=466205 $Y=492465 $D=0
M9 4 37 243 4 N L=1.8e-07 W=5.7e-07 $X=466925 $Y=492465 $D=0
M10 243 37 4 4 N L=1.8e-07 W=5.7e-07 $X=467645 $Y=492465 $D=0
M11 4 37 243 4 N L=1.8e-07 W=5.7e-07 $X=468365 $Y=492465 $D=0
M12 243 37 4 4 N L=1.8e-07 W=5.7e-07 $X=469085 $Y=492465 $D=0
M13 4 37 243 4 N L=1.8e-07 W=5.7e-07 $X=469805 $Y=492465 $D=0
M14 243 253 4 4 N L=1.8e-07 W=5.7e-07 $X=470525 $Y=492465 $D=0
M15 4 253 243 4 N L=1.8e-07 W=5.7e-07 $X=471245 $Y=492465 $D=0
M16 243 253 4 4 N L=1.8e-07 W=5.7e-07 $X=471965 $Y=492465 $D=0
M17 4 253 243 4 N L=1.8e-07 W=5.7e-07 $X=472685 $Y=492465 $D=0
M18 243 253 4 4 N L=1.8e-07 W=5.7e-07 $X=473405 $Y=492465 $D=0
M19 4 253 243 4 N L=1.8e-07 W=5.7e-07 $X=474125 $Y=492465 $D=0
M20 243 253 4 4 N L=1.8e-07 W=5.7e-07 $X=474845 $Y=492465 $D=0
M21 555 26 4 4 N L=1.8e-07 W=1e-06 $X=478740 $Y=584855 $D=0
M22 556 60 555 4 N L=1.8e-07 W=1e-06 $X=479515 $Y=584855 $D=0
M23 265 31 556 4 N L=1.8e-07 W=1e-06 $X=480285 $Y=584855 $D=0
M24 557 31 265 4 N L=1.8e-07 W=1e-06 $X=481005 $Y=584855 $D=0
M25 558 60 557 4 N L=1.8e-07 W=1e-06 $X=481685 $Y=584855 $D=0
M26 4 26 558 4 N L=1.8e-07 W=1e-06 $X=482365 $Y=584855 $D=0
M27 24 265 4 4 N L=1.8e-07 W=1e-06 $X=483325 $Y=584855 $D=0
M28 4 265 24 4 N L=1.8e-07 W=1e-06 $X=484045 $Y=584855 $D=0
M29 24 265 4 4 N L=1.8e-07 W=1e-06 $X=484905 $Y=584855 $D=0
M30 4 265 24 4 N L=1.8e-07 W=1e-06 $X=485625 $Y=584855 $D=0
M31 4 297 292 4 N L=1.8e-07 W=5e-07 $X=510660 $Y=563140 $D=0
M32 297 296 4 4 N L=1.8e-07 W=5e-07 $X=511380 $Y=563140 $D=0
M33 559 286 297 4 N L=1.8e-07 W=5e-07 $X=512100 $Y=563140 $D=0
M34 4 260 559 4 N L=1.8e-07 W=5e-07 $X=512600 $Y=563140 $D=0
M35 393 376 4 4 N L=1.8e-07 W=1e-06 $X=581220 $Y=490775 $D=0
M36 4 384 393 4 N L=1.8e-07 W=1e-06 $X=581940 $Y=490775 $D=0
M37 396 393 4 4 N L=1.8e-07 W=1e-06 $X=582750 $Y=490775 $D=0
M38 560 384 396 4 N L=1.8e-07 W=1e-06 $X=583555 $Y=490775 $D=0
M39 4 376 560 4 N L=1.8e-07 W=1e-06 $X=584280 $Y=490775 $D=0
M40 245 41 1 1 P L=1.8e-07 W=1.36e-06 $X=460445 $Y=494335 $D=16
M41 1 41 245 1 P L=1.8e-07 W=1.6e-06 $X=461165 $Y=494095 $D=16
M42 245 41 1 1 P L=1.8e-07 W=1.6e-06 $X=461885 $Y=494095 $D=16
M43 1 41 245 1 P L=1.8e-07 W=1.6e-06 $X=462605 $Y=494095 $D=16
M44 245 41 1 1 P L=1.8e-07 W=1.6e-06 $X=463325 $Y=494095 $D=16
M45 1 41 245 1 P L=1.8e-07 W=1.6e-06 $X=464045 $Y=494095 $D=16
M46 245 41 1 1 P L=1.8e-07 W=1.6e-06 $X=464765 $Y=494095 $D=16
M47 250 37 245 1 P L=1.8e-07 W=1.6e-06 $X=465485 $Y=494095 $D=16
M48 245 37 250 1 P L=1.8e-07 W=1.6e-06 $X=466205 $Y=494095 $D=16
M49 250 37 245 1 P L=1.8e-07 W=1.6e-06 $X=466925 $Y=494095 $D=16
M50 245 37 250 1 P L=1.8e-07 W=1.6e-06 $X=467645 $Y=494095 $D=16
M51 250 37 245 1 P L=1.8e-07 W=1.6e-06 $X=468365 $Y=494095 $D=16
M52 245 37 250 1 P L=1.8e-07 W=1.6e-06 $X=469085 $Y=494095 $D=16
M53 250 37 245 1 P L=1.8e-07 W=1.6e-06 $X=469805 $Y=494095 $D=16
M54 243 253 250 1 P L=1.8e-07 W=1.6e-06 $X=470525 $Y=494095 $D=16
M55 250 253 243 1 P L=1.8e-07 W=1.6e-06 $X=471245 $Y=494095 $D=16
M56 243 253 250 1 P L=1.8e-07 W=1.6e-06 $X=471965 $Y=494095 $D=16
M57 250 253 243 1 P L=1.8e-07 W=1.6e-06 $X=472685 $Y=494095 $D=16
M58 243 253 250 1 P L=1.8e-07 W=1.6e-06 $X=473405 $Y=494095 $D=16
M59 250 253 243 1 P L=1.8e-07 W=1.6e-06 $X=474125 $Y=494095 $D=16
M60 243 253 250 1 P L=1.8e-07 W=1.36e-06 $X=474845 $Y=494335 $D=16
M61 265 26 1 1 P L=1.8e-07 W=1.37e-06 $X=478740 $Y=582625 $D=16
M62 1 60 265 1 P L=1.8e-07 W=1.37e-06 $X=479460 $Y=582625 $D=16
M63 265 31 1 1 P L=1.8e-07 W=1.37e-06 $X=480285 $Y=582625 $D=16
M64 1 31 265 1 P L=1.8e-07 W=1.37e-06 $X=481005 $Y=582625 $D=16
M65 265 60 1 1 P L=1.8e-07 W=1.37e-06 $X=481805 $Y=582625 $D=16
M66 1 26 265 1 P L=1.8e-07 W=1.37e-06 $X=482525 $Y=582625 $D=16
M67 24 265 1 1 P L=1.8e-07 W=1.37e-06 $X=483325 $Y=582625 $D=16
M68 1 265 24 1 P L=1.8e-07 W=1.37e-06 $X=484045 $Y=582625 $D=16
M69 24 265 1 1 P L=1.8e-07 W=1.37e-06 $X=484905 $Y=582625 $D=16
M70 1 265 24 1 P L=1.8e-07 W=1.37e-06 $X=485625 $Y=582625 $D=16
M71 1 297 292 1 P L=1.8e-07 W=6.85e-07 $X=510660 $Y=565235 $D=16
M72 561 296 1 1 P L=1.8e-07 W=6.85e-07 $X=511380 $Y=565235 $D=16
M73 297 286 561 1 P L=1.8e-07 W=6.85e-07 $X=512010 $Y=565235 $D=16
M74 561 260 297 1 P L=1.8e-07 W=6.85e-07 $X=512730 $Y=565235 $D=16
M75 562 376 393 1 P L=1.8e-07 W=1.37e-06 $X=581220 $Y=488545 $D=16
M76 1 384 562 1 P L=1.8e-07 W=1.37e-06 $X=581930 $Y=488545 $D=16
M77 394 393 1 1 P L=1.8e-07 W=1.37e-06 $X=582750 $Y=488545 $D=16
M78 396 384 394 1 P L=1.8e-07 W=1.37e-06 $X=583555 $Y=488545 $D=16
M79 394 376 396 1 P L=1.8e-07 W=1.37e-06 $X=584280 $Y=488545 $D=16
X273 1 4 DCAPBWP7T $T=458520 523480 1 0 $X=458230 $Y=519270
X274 1 4 DCAPBWP7T $T=468040 515640 0 0 $X=467750 $Y=515405
X275 1 4 DCAPBWP7T $T=468600 562680 1 0 $X=468310 $Y=558470
X276 1 4 DCAPBWP7T $T=475880 531320 0 0 $X=475590 $Y=531085
X277 1 4 DCAPBWP7T $T=480360 492120 0 0 $X=480070 $Y=491885
X278 1 4 DCAPBWP7T $T=481480 515640 1 0 $X=481190 $Y=511430
X279 1 4 DCAPBWP7T $T=481480 562680 1 0 $X=481190 $Y=558470
X280 1 4 DCAPBWP7T $T=482040 570520 0 0 $X=481750 $Y=570285
X281 1 4 DCAPBWP7T $T=489320 539160 0 0 $X=489030 $Y=538925
X282 1 4 DCAPBWP7T $T=489320 578360 1 0 $X=489030 $Y=574150
X283 1 4 DCAPBWP7T $T=494360 515640 0 0 $X=494070 $Y=515405
X284 1 4 DCAPBWP7T $T=498840 586200 0 0 $X=498550 $Y=585965
X285 1 4 DCAPBWP7T $T=506120 499960 1 0 $X=505830 $Y=495750
X286 1 4 DCAPBWP7T $T=507240 523480 1 0 $X=506950 $Y=519270
X287 1 4 DCAPBWP7T $T=512280 554840 1 0 $X=511990 $Y=550630
X288 1 4 DCAPBWP7T $T=513960 515640 1 0 $X=513670 $Y=511430
X289 1 4 DCAPBWP7T $T=514520 492120 0 0 $X=514230 $Y=491885
X290 1 4 DCAPBWP7T $T=514520 531320 0 0 $X=514230 $Y=531085
X291 1 4 DCAPBWP7T $T=524600 562680 1 0 $X=524310 $Y=558470
X292 1 4 DCAPBWP7T $T=531320 523480 1 0 $X=531030 $Y=519270
X293 1 4 DCAPBWP7T $T=531320 531320 0 0 $X=531030 $Y=531085
X294 1 4 DCAPBWP7T $T=531320 578360 1 0 $X=531030 $Y=574150
X295 1 4 DCAPBWP7T $T=540840 539160 0 0 $X=540550 $Y=538925
X296 1 4 DCAPBWP7T $T=543080 492120 1 0 $X=542790 $Y=487910
X297 1 4 DCAPBWP7T $T=552040 499960 1 0 $X=551750 $Y=495750
X298 1 4 DCAPBWP7T $T=583400 484280 0 0 $X=583110 $Y=484045
X299 1 4 DCAPBWP7T $T=585080 578360 0 0 $X=584790 $Y=578125
X300 1 4 DCAPBWP7T $T=601320 539160 0 0 $X=601030 $Y=538925
X301 1 4 DCAPBWP7T $T=605240 594040 1 0 $X=604950 $Y=589830
X302 1 4 DCAPBWP7T $T=608040 523480 0 0 $X=607750 $Y=523245
X303 1 4 DCAPBWP7T $T=608040 539160 0 0 $X=607750 $Y=538925
X304 1 4 DCAPBWP7T $T=615320 547000 1 0 $X=615030 $Y=542790
X305 1 4 DCAPBWP7T $T=618120 492120 0 0 $X=617830 $Y=491885
X306 1 4 DCAPBWP7T $T=618120 594040 1 0 $X=617830 $Y=589830
X307 1 4 DCAPBWP7T $T=620360 507800 1 0 $X=620070 $Y=503590
X308 1 4 DCAPBWP7T $T=622600 523480 1 0 $X=622310 $Y=519270
X309 1 4 DCAPBWP7T $T=631560 492120 1 0 $X=631270 $Y=487910
X310 1 4 DCAPBWP7T $T=636040 515640 1 0 $X=635750 $Y=511430
X311 1 4 DCAPBWP7T $T=646120 539160 1 0 $X=645830 $Y=534950
X312 1 4 DCAPBWP7T $T=647800 515640 0 0 $X=647510 $Y=515405
X313 1 4 DCAPBWP7T $T=647800 531320 0 0 $X=647510 $Y=531085
X314 1 4 DCAPBWP7T $T=650040 523480 0 0 $X=649750 $Y=523245
X315 1 4 DCAPBWP7T $T=657320 492120 0 0 $X=657030 $Y=491885
X316 1 4 DCAPBWP7T $T=657320 507800 1 0 $X=657030 $Y=503590
X317 1 4 DCAPBWP7T $T=657320 515640 1 0 $X=657030 $Y=511430
X318 1 4 DCAPBWP7T $T=657320 539160 1 0 $X=657030 $Y=534950
X319 1 4 DCAPBWP7T $T=657320 547000 0 0 $X=657030 $Y=546765
X320 1 4 DCAPBWP7T $T=657320 554840 1 0 $X=657030 $Y=550630
X321 1 4 DCAPBWP7T $T=669640 515640 1 0 $X=669350 $Y=511430
X322 1 4 DCAPBWP7T $T=680280 531320 0 0 $X=679990 $Y=531085
X323 1 4 DCAPBWP7T $T=684200 499960 0 0 $X=683910 $Y=499725
X324 1 4 DCAPBWP7T $T=684760 523480 1 0 $X=684470 $Y=519270
X325 1 4 DCAPBWP7T $T=687000 594040 0 0 $X=686710 $Y=593805
X326 1 4 DCAPBWP7T $T=691480 539160 0 0 $X=691190 $Y=538925
X327 1 4 DCAPBWP7T $T=699320 484280 0 0 $X=699030 $Y=484045
X328 1 4 DCAPBWP7T $T=699320 499960 1 0 $X=699030 $Y=495750
X329 1 4 DCAPBWP7T $T=699320 515640 1 0 $X=699030 $Y=511430
X330 1 4 DCAPBWP7T $T=699320 531320 1 0 $X=699030 $Y=527110
X331 1 4 DCAPBWP7T $T=699320 570520 0 0 $X=699030 $Y=570285
X332 1 4 DCAPBWP7T $T=699320 586200 0 0 $X=699030 $Y=585965
X333 1 4 DCAPBWP7T $T=713320 586200 1 0 $X=713030 $Y=581990
X334 1 4 DCAPBWP7T $T=717800 554840 1 0 $X=717510 $Y=550630
X335 1 4 DCAPBWP7T $T=722280 594040 1 0 $X=721990 $Y=589830
X336 1 4 DCAPBWP7T $T=722840 484280 0 0 $X=722550 $Y=484045
X337 1 4 DCAPBWP7T $T=733480 531320 1 0 $X=733190 $Y=527110
X338 1 4 DCAPBWP7T $T=734600 554840 0 0 $X=734310 $Y=554605
X339 1 4 DCAPBWP7T $T=741320 499960 0 0 $X=741030 $Y=499725
X340 1 4 DCAPBWP7T $T=741320 578360 1 0 $X=741030 $Y=574150
X341 1 4 DCAPBWP7T $T=741320 586200 1 0 $X=741030 $Y=581990
X342 4 1 DCAP8BWP7T $T=450120 594040 0 0 $X=449830 $Y=593805
X343 4 1 DCAP8BWP7T $T=463560 499960 1 0 $X=463270 $Y=495750
X344 4 1 DCAP8BWP7T $T=475880 492120 0 0 $X=475590 $Y=491885
X345 4 1 DCAP8BWP7T $T=485960 523480 0 0 $X=485670 $Y=523245
X346 4 1 DCAP8BWP7T $T=485960 531320 1 0 $X=485670 $Y=527110
X347 4 1 DCAP8BWP7T $T=492120 570520 0 0 $X=491830 $Y=570285
X348 4 1 DCAP8BWP7T $T=501080 562680 0 0 $X=500790 $Y=562445
X349 4 1 DCAP8BWP7T $T=502200 492120 1 0 $X=501910 $Y=487910
X350 4 1 DCAP8BWP7T $T=503320 547000 0 0 $X=503030 $Y=546765
X351 4 1 DCAP8BWP7T $T=507240 523480 0 0 $X=506950 $Y=523245
X352 4 1 DCAP8BWP7T $T=510040 492120 0 0 $X=509750 $Y=491885
X353 4 1 DCAP8BWP7T $T=510040 594040 1 0 $X=509750 $Y=589830
X354 4 1 DCAP8BWP7T $T=525720 499960 1 0 $X=525430 $Y=495750
X355 4 1 DCAP8BWP7T $T=526840 531320 0 0 $X=526550 $Y=531085
X356 4 1 DCAP8BWP7T $T=527960 492120 1 0 $X=527670 $Y=487910
X357 4 1 DCAP8BWP7T $T=543080 523480 1 0 $X=542790 $Y=519270
X358 4 1 DCAP8BWP7T $T=547560 499960 1 0 $X=547270 $Y=495750
X359 4 1 DCAP8BWP7T $T=569960 515640 0 0 $X=569670 $Y=515405
X360 4 1 DCAP8BWP7T $T=569960 523480 1 0 $X=569670 $Y=519270
X361 4 1 DCAP8BWP7T $T=569960 586200 1 0 $X=569670 $Y=581990
X362 4 1 DCAP8BWP7T $T=594040 554840 1 0 $X=593750 $Y=550630
X363 4 1 DCAP8BWP7T $T=611960 554840 1 0 $X=611670 $Y=550630
X364 4 1 DCAP8BWP7T $T=611960 570520 1 0 $X=611670 $Y=566310
X365 4 1 DCAP8BWP7T $T=618120 523480 1 0 $X=617830 $Y=519270
X366 4 1 DCAP8BWP7T $T=636040 547000 1 0 $X=635750 $Y=542790
X367 4 1 DCAP8BWP7T $T=641080 570520 0 0 $X=640790 $Y=570285
X368 4 1 DCAP8BWP7T $T=641640 539160 1 0 $X=641350 $Y=534950
X369 4 1 DCAP8BWP7T $T=652840 492120 0 0 $X=652550 $Y=491885
X370 4 1 DCAP8BWP7T $T=653960 499960 1 0 $X=653670 $Y=495750
X371 4 1 DCAP8BWP7T $T=660120 499960 0 0 $X=659830 $Y=499725
X372 4 1 DCAP8BWP7T $T=660120 562680 0 0 $X=659830 $Y=562445
X373 4 1 DCAP8BWP7T $T=669080 523480 0 0 $X=668790 $Y=523245
X374 4 1 DCAP8BWP7T $T=684760 578360 1 0 $X=684470 $Y=574150
X375 4 1 DCAP8BWP7T $T=686440 507800 0 0 $X=686150 $Y=507565
X376 4 1 DCAP8BWP7T $T=687000 539160 0 0 $X=686710 $Y=538925
X377 4 1 DCAP8BWP7T $T=687000 586200 0 0 $X=686710 $Y=585965
X378 4 1 DCAP8BWP7T $T=694840 586200 0 0 $X=694550 $Y=585965
X379 4 1 DCAP8BWP7T $T=702120 539160 0 0 $X=701830 $Y=538925
X380 4 1 DCAP8BWP7T $T=718360 484280 0 0 $X=718070 $Y=484045
X381 4 1 DCAP8BWP7T $T=719480 570520 1 0 $X=719190 $Y=566310
X382 4 1 DCAP8BWP7T $T=720040 578360 1 0 $X=719750 $Y=574150
X383 4 1 DCAP8BWP7T $T=723400 492120 0 0 $X=723110 $Y=491885
X384 4 1 DCAP8BWP7T $T=730120 554840 0 0 $X=729830 $Y=554605
X385 4 1 DCAP8BWP7T $T=736840 578360 1 0 $X=736550 $Y=574150
X386 4 1 DCAP8BWP7T $T=737960 594040 0 0 $X=737670 $Y=593805
X387 4 1 DCAP4BWP7T $T=459080 507800 1 0 $X=458790 $Y=503590
X388 4 1 DCAP4BWP7T $T=477000 547000 1 0 $X=476710 $Y=542790
X389 4 1 DCAP4BWP7T $T=487080 578360 1 0 $X=486790 $Y=574150
X390 4 1 DCAP4BWP7T $T=488200 499960 1 0 $X=487910 $Y=495750
X391 4 1 DCAP4BWP7T $T=488760 547000 0 0 $X=488470 $Y=546765
X392 4 1 DCAP4BWP7T $T=488760 562680 0 0 $X=488470 $Y=562445
X393 4 1 DCAP4BWP7T $T=492120 499960 0 0 $X=491830 $Y=499725
X394 4 1 DCAP4BWP7T $T=492120 515640 0 0 $X=491830 $Y=515405
X395 4 1 DCAP4BWP7T $T=492120 523480 1 0 $X=491830 $Y=519270
X396 4 1 DCAP4BWP7T $T=503880 499960 1 0 $X=503590 $Y=495750
X397 4 1 DCAP4BWP7T $T=503880 539160 1 0 $X=503590 $Y=534950
X398 4 1 DCAP4BWP7T $T=512280 531320 0 0 $X=511990 $Y=531085
X399 4 1 DCAP4BWP7T $T=520680 499960 1 0 $X=520390 $Y=495750
X400 4 1 DCAP4BWP7T $T=524040 484280 0 0 $X=523750 $Y=484045
X401 4 1 DCAP4BWP7T $T=530200 539160 0 0 $X=529910 $Y=538925
X402 4 1 DCAP4BWP7T $T=530760 507800 0 0 $X=530470 $Y=507565
X403 4 1 DCAP4BWP7T $T=530760 547000 1 0 $X=530470 $Y=542790
X404 4 1 DCAP4BWP7T $T=530760 547000 0 0 $X=530470 $Y=546765
X405 4 1 DCAP4BWP7T $T=534120 515640 0 0 $X=533830 $Y=515405
X406 4 1 DCAP4BWP7T $T=534120 531320 1 0 $X=533830 $Y=527110
X407 4 1 DCAP4BWP7T $T=552040 547000 0 0 $X=551750 $Y=546765
X408 4 1 DCAP4BWP7T $T=572200 547000 1 0 $X=571910 $Y=542790
X409 4 1 DCAP4BWP7T $T=572200 594040 0 0 $X=571910 $Y=593805
X410 4 1 DCAP4BWP7T $T=572760 562680 1 0 $X=572470 $Y=558470
X411 4 1 DCAP4BWP7T $T=592360 554840 0 0 $X=592070 $Y=554605
X412 4 1 DCAP4BWP7T $T=594040 523480 1 0 $X=593750 $Y=519270
X413 4 1 DCAP4BWP7T $T=605800 523480 0 0 $X=605510 $Y=523245
X414 4 1 DCAP4BWP7T $T=614200 539160 1 0 $X=613910 $Y=534950
X415 4 1 DCAP4BWP7T $T=614200 547000 0 0 $X=613910 $Y=546765
X416 4 1 DCAP4BWP7T $T=618120 507800 1 0 $X=617830 $Y=503590
X417 4 1 DCAP4BWP7T $T=637160 531320 0 0 $X=636870 $Y=531085
X418 4 1 DCAP4BWP7T $T=656200 484280 0 0 $X=655910 $Y=484045
X419 4 1 DCAP4BWP7T $T=656200 586200 0 0 $X=655910 $Y=585965
X420 4 1 DCAP4BWP7T $T=660120 499960 1 0 $X=659830 $Y=495750
X421 4 1 DCAP4BWP7T $T=660120 586200 0 0 $X=659830 $Y=585965
X422 4 1 DCAP4BWP7T $T=671880 578360 1 0 $X=671590 $Y=574150
X423 4 1 DCAP4BWP7T $T=678040 531320 0 0 $X=677750 $Y=531085
X424 4 1 DCAP4BWP7T $T=682520 523480 1 0 $X=682230 $Y=519270
X425 4 1 DCAP4BWP7T $T=697080 484280 0 0 $X=696790 $Y=484045
X426 4 1 DCAP4BWP7T $T=698200 547000 0 0 $X=697910 $Y=546765
X427 4 1 DCAP4BWP7T $T=698200 554840 0 0 $X=697910 $Y=554605
X428 4 1 DCAP4BWP7T $T=698760 523480 1 0 $X=698470 $Y=519270
X429 4 1 DCAP4BWP7T $T=698760 594040 1 0 $X=698470 $Y=589830
X430 4 1 DCAP4BWP7T $T=711080 586200 1 0 $X=710790 $Y=581990
X431 4 1 DCAP4BWP7T $T=715560 554840 1 0 $X=715270 $Y=550630
X432 4 1 DCAP4BWP7T $T=721160 523480 0 0 $X=720870 $Y=523245
X433 4 1 DCAP4BWP7T $T=731240 531320 1 0 $X=730950 $Y=527110
X434 4 1 DCAP4BWP7T $T=733480 515640 1 0 $X=733190 $Y=511430
X435 4 1 DCAP4BWP7T $T=740760 515640 0 0 $X=740470 $Y=515405
X436 4 1 DCAP4BWP7T $T=740760 554840 1 0 $X=740470 $Y=550630
X437 4 1 ICV_40 $T=450120 562680 1 0 $X=449830 $Y=558470
X438 4 1 ICV_40 $T=461880 562680 1 0 $X=461590 $Y=558470
X439 4 1 ICV_40 $T=468040 531320 1 0 $X=467750 $Y=527110
X440 4 1 ICV_40 $T=468040 570520 1 0 $X=467750 $Y=566310
X441 4 1 ICV_40 $T=482600 539160 0 0 $X=482310 $Y=538925
X442 4 1 ICV_40 $T=484280 499960 0 0 $X=483990 $Y=499725
X443 4 1 ICV_40 $T=484280 547000 1 0 $X=483990 $Y=542790
X444 4 1 ICV_40 $T=492120 562680 0 0 $X=491830 $Y=562445
X445 4 1 ICV_40 $T=492120 586200 0 0 $X=491830 $Y=585965
X446 4 1 ICV_40 $T=501640 499960 0 0 $X=501350 $Y=499725
X447 4 1 ICV_40 $T=511160 586200 0 0 $X=510870 $Y=585965
X448 4 1 ICV_40 $T=517880 562680 1 0 $X=517590 $Y=558470
X449 4 1 ICV_40 $T=519000 586200 1 0 $X=518710 $Y=581990
X450 4 1 ICV_40 $T=525720 594040 1 0 $X=525430 $Y=589830
X451 4 1 ICV_40 $T=526280 515640 0 0 $X=525990 $Y=515405
X452 4 1 ICV_40 $T=526280 539160 1 0 $X=525990 $Y=534950
X453 4 1 ICV_40 $T=526280 570520 1 0 $X=525990 $Y=566310
X454 4 1 ICV_40 $T=534120 539160 0 0 $X=533830 $Y=538925
X455 4 1 ICV_40 $T=585080 594040 1 0 $X=584790 $Y=589830
X456 4 1 ICV_40 $T=608600 547000 1 0 $X=608310 $Y=542790
X457 4 1 ICV_40 $T=609720 570520 0 0 $X=609430 $Y=570285
X458 4 1 ICV_40 $T=610280 531320 0 0 $X=609990 $Y=531085
X459 4 1 ICV_40 $T=618120 515640 1 0 $X=617830 $Y=511430
X460 4 1 ICV_40 $T=623720 492120 0 0 $X=623430 $Y=491885
X461 4 1 ICV_40 $T=623720 507800 1 0 $X=623430 $Y=503590
X462 4 1 ICV_40 $T=635480 492120 0 0 $X=635190 $Y=491885
X463 4 1 ICV_40 $T=642200 507800 0 0 $X=641910 $Y=507565
X464 4 1 ICV_40 $T=650600 539160 1 0 $X=650310 $Y=534950
X465 4 1 ICV_40 $T=650600 547000 0 0 $X=650310 $Y=546765
X466 4 1 ICV_40 $T=651720 531320 0 0 $X=651430 $Y=531085
X467 4 1 ICV_40 $T=652280 507800 0 0 $X=651990 $Y=507565
X468 4 1 ICV_40 $T=652280 515640 0 0 $X=651990 $Y=515405
X469 4 1 ICV_40 $T=660120 484280 0 0 $X=659830 $Y=484045
X470 4 1 ICV_40 $T=660120 523480 0 0 $X=659830 $Y=523245
X471 4 1 ICV_40 $T=660120 547000 0 0 $X=659830 $Y=546765
X472 4 1 ICV_40 $T=660120 594040 1 0 $X=659830 $Y=589830
X473 4 1 ICV_40 $T=669080 554840 0 0 $X=668790 $Y=554605
X474 4 1 ICV_40 $T=677480 499960 0 0 $X=677190 $Y=499725
X475 4 1 ICV_40 $T=685320 554840 1 0 $X=685030 $Y=550630
X476 4 1 ICV_40 $T=686440 523480 0 0 $X=686150 $Y=523245
X477 4 1 ICV_40 $T=692600 515640 1 0 $X=692310 $Y=511430
X478 4 1 ICV_40 $T=693720 507800 0 0 $X=693430 $Y=507565
X479 4 1 ICV_40 $T=694280 578360 1 0 $X=693990 $Y=574150
X480 4 1 ICV_40 $T=702120 523480 0 0 $X=701830 $Y=523245
X481 4 1 ICV_40 $T=711080 499960 1 0 $X=710790 $Y=495750
X482 4 1 ICV_40 $T=727320 484280 0 0 $X=727030 $Y=484045
X483 4 1 ICV_40 $T=734600 586200 1 0 $X=734310 $Y=581990
X484 4 1 ICV_40 $T=736280 492120 1 0 $X=735990 $Y=487910
X485 4 1 ICV_40 $T=736280 507800 0 0 $X=735990 $Y=507565
X486 4 1 ICV_40 $T=736280 523480 0 0 $X=735990 $Y=523245
X487 4 1 ICV_40 $T=736280 570520 1 0 $X=735990 $Y=566310
X488 231 1 232 229 4 NR2D1BWP7T $T=458520 523480 0 180 $X=455990 $Y=519270
X489 240 1 241 48 4 NR2D1BWP7T $T=464120 547000 1 0 $X=463830 $Y=542790
X490 244 1 242 23 4 NR2D1BWP7T $T=469160 531320 1 180 $X=466630 $Y=531085
X491 259 1 256 23 4 NR2D1BWP7T $T=481480 547000 0 180 $X=478950 $Y=542790
X492 67 1 268 23 4 NR2D1BWP7T $T=485400 515640 0 180 $X=482870 $Y=511430
X493 68 1 246 23 4 NR2D1BWP7T $T=485400 562680 0 180 $X=482870 $Y=558470
X494 74 1 254 71 4 NR2D1BWP7T $T=494920 539160 0 180 $X=492390 $Y=534950
X495 74 1 273 23 4 NR2D1BWP7T $T=496040 547000 0 180 $X=493510 $Y=542790
X496 48 1 233 23 4 NR2D1BWP7T $T=501080 562680 1 180 $X=498550 $Y=562445
X497 33 1 78 253 4 NR2D1BWP7T $T=503880 499960 0 180 $X=501350 $Y=495750
X498 74 1 283 259 4 NR2D1BWP7T $T=502200 578360 1 0 $X=501910 $Y=574150
X499 71 1 299 240 4 NR2D1BWP7T $T=506120 539160 1 0 $X=505830 $Y=534950
X500 74 1 290 249 4 NR2D1BWP7T $T=507800 554840 1 0 $X=507510 $Y=550630
X501 19 1 294 295 4 NR2D1BWP7T $T=509480 515640 1 0 $X=509190 $Y=511430
X502 240 1 300 23 4 NR2D1BWP7T $T=513960 562680 0 0 $X=513670 $Y=562445
X503 240 1 301 249 4 NR2D1BWP7T $T=513960 578360 1 0 $X=513670 $Y=574150
X504 87 1 287 88 4 NR2D1BWP7T $T=516200 492120 0 0 $X=515910 $Y=491885
X505 88 1 305 65 4 NR2D1BWP7T $T=519560 484280 1 180 $X=517030 $Y=484045
X506 71 1 312 99 4 NR2D1BWP7T $T=524040 570520 1 0 $X=523750 $Y=566310
X507 71 1 314 101 4 NR2D1BWP7T $T=524600 578360 1 0 $X=524310 $Y=574150
X508 87 1 316 100 4 NR2D1BWP7T $T=525720 492120 1 0 $X=525430 $Y=487910
X509 100 1 320 65 4 NR2D1BWP7T $T=526280 484280 0 0 $X=525990 $Y=484045
X510 71 1 318 104 4 NR2D1BWP7T $T=526280 554840 0 0 $X=525990 $Y=554605
X511 259 1 319 240 4 NR2D1BWP7T $T=526280 562680 1 0 $X=525990 $Y=558470
X512 240 1 322 68 4 NR2D1BWP7T $T=526280 578360 0 0 $X=525990 $Y=578125
X513 249 1 103 99 4 NR2D1BWP7T $T=526280 586200 1 0 $X=525990 $Y=581990
X514 104 1 328 48 4 NR2D1BWP7T $T=536360 554840 0 0 $X=536070 $Y=554605
X515 100 1 330 23 4 NR2D1BWP7T $T=536920 484280 0 0 $X=536630 $Y=484045
X516 71 1 344 108 4 NR2D1BWP7T $T=550360 570520 0 0 $X=550070 $Y=570285
X517 99 1 351 110 4 NR2D1BWP7T $T=552600 570520 0 0 $X=552310 $Y=570285
X518 74 1 354 244 4 NR2D1BWP7T $T=554840 570520 0 0 $X=554550 $Y=570285
X519 87 1 121 392 4 NR2D1BWP7T $T=576680 484280 0 0 $X=576390 $Y=484045
X520 104 1 122 110 4 NR2D1BWP7T $T=576680 578360 1 0 $X=576390 $Y=574150
X521 249 1 390 108 4 NR2D1BWP7T $T=578920 578360 1 0 $X=578630 $Y=574150
X522 88 1 370 125 4 NR2D1BWP7T $T=585080 484280 0 0 $X=584790 $Y=484045
X523 88 1 386 23 4 NR2D1BWP7T $T=603000 515640 0 0 $X=602710 $Y=515405
X524 392 1 371 23 4 NR2D1BWP7T $T=608040 515640 1 180 $X=605510 $Y=515405
X525 142 1 429 65 4 NR2D1BWP7T $T=606920 484280 0 0 $X=606630 $Y=484045
X526 143 1 424 65 4 NR2D1BWP7T $T=609160 492120 0 180 $X=606630 $Y=487910
X527 240 1 420 110 4 NR2D1BWP7T $T=609160 594040 0 180 $X=606630 $Y=589830
X528 422 1 432 149 4 NR2D1BWP7T $T=609160 515640 0 0 $X=608870 $Y=515405
X529 104 1 409 68 4 NR2D1BWP7T $T=610280 562680 0 0 $X=609990 $Y=562445
X530 143 1 412 23 4 NR2D1BWP7T $T=620920 515640 1 180 $X=618390 $Y=515405
X531 104 1 348 249 4 NR2D1BWP7T $T=621480 578360 0 180 $X=618950 $Y=574150
X532 101 1 436 48 4 NR2D1BWP7T $T=620920 578360 0 0 $X=620630 $Y=578125
X533 157 1 402 23 4 NR2D1BWP7T $T=626520 523480 0 180 $X=623990 $Y=519270
X534 142 1 403 23 4 NR2D1BWP7T $T=647800 523480 0 0 $X=647510 $Y=523245
X535 1 4 DCAP64BWP7T $T=452920 562680 0 0 $X=452630 $Y=562445
X536 1 4 DCAP64BWP7T $T=581160 578360 1 0 $X=580870 $Y=574150
X537 1 4 DCAP64BWP7T $T=664040 570520 1 0 $X=663750 $Y=566310
X577 4 1 ICV_47 $T=450120 484280 0 0 $X=449830 $Y=484045
X578 4 1 ICV_47 $T=450120 539160 1 0 $X=449830 $Y=534950
X579 4 1 ICV_47 $T=450120 554840 1 0 $X=449830 $Y=550630
X580 4 1 ICV_47 $T=450120 578360 0 0 $X=449830 $Y=578125
X581 4 1 ICV_47 $T=450120 586200 0 0 $X=449830 $Y=585965
X582 4 1 ICV_47 $T=534120 492120 0 0 $X=533830 $Y=491885
X583 4 1 ICV_47 $T=534120 507800 1 0 $X=533830 $Y=503590
X584 4 1 ICV_47 $T=534120 531320 0 0 $X=533830 $Y=531085
X585 4 1 ICV_47 $T=534120 539160 1 0 $X=533830 $Y=534950
X586 4 1 ICV_47 $T=534120 554840 1 0 $X=533830 $Y=550630
X587 4 1 ICV_47 $T=534120 578360 0 0 $X=533830 $Y=578125
X588 4 1 ICV_47 $T=576120 492120 0 0 $X=575830 $Y=491885
X589 4 1 ICV_47 $T=576120 586200 1 0 $X=575830 $Y=581990
X590 4 1 ICV_47 $T=618120 499960 0 0 $X=617830 $Y=499725
X591 4 1 ICV_47 $T=618120 539160 0 0 $X=617830 $Y=538925
X592 4 1 ICV_47 $T=618120 554840 0 0 $X=617830 $Y=554605
X593 4 1 ICV_47 $T=618120 570520 1 0 $X=617830 $Y=566310
X594 4 1 ICV_47 $T=618120 586200 1 0 $X=617830 $Y=581990
X595 4 1 ICV_47 $T=618120 594040 0 0 $X=617830 $Y=593805
X596 4 1 ICV_47 $T=660120 492120 0 0 $X=659830 $Y=491885
X597 4 1 ICV_47 $T=660120 507800 1 0 $X=659830 $Y=503590
X598 4 1 ICV_47 $T=660120 547000 1 0 $X=659830 $Y=542790
X599 4 1 ICV_47 $T=660120 586200 1 0 $X=659830 $Y=581990
X600 4 1 ICV_47 $T=702120 586200 0 0 $X=701830 $Y=585965
X601 1 4 DCAP32BWP7T $T=450120 492120 1 0 $X=449830 $Y=487910
X602 1 4 DCAP32BWP7T $T=450120 499960 0 0 $X=449830 $Y=499725
X603 1 4 DCAP32BWP7T $T=450120 515640 1 0 $X=449830 $Y=511430
X604 1 4 DCAP32BWP7T $T=450120 515640 0 0 $X=449830 $Y=515405
X605 1 4 DCAP32BWP7T $T=450120 531320 1 0 $X=449830 $Y=527110
X606 1 4 DCAP32BWP7T $T=450120 570520 1 0 $X=449830 $Y=566310
X607 1 4 DCAP32BWP7T $T=492120 492120 0 0 $X=491830 $Y=491885
X608 1 4 DCAP32BWP7T $T=496040 547000 1 0 $X=495750 $Y=542790
X609 1 4 DCAP32BWP7T $T=507240 531320 1 0 $X=506950 $Y=527110
X610 1 4 DCAP32BWP7T $T=534120 547000 0 0 $X=533830 $Y=546765
X611 1 4 DCAP32BWP7T $T=534120 562680 0 0 $X=533830 $Y=562445
X612 1 4 DCAP32BWP7T $T=534120 578360 1 0 $X=533830 $Y=574150
X613 1 4 DCAP32BWP7T $T=534120 594040 1 0 $X=533830 $Y=589830
X614 1 4 DCAP32BWP7T $T=539160 515640 0 0 $X=538870 $Y=515405
X615 1 4 DCAP32BWP7T $T=551480 554840 0 0 $X=551190 $Y=554605
X616 1 4 DCAP32BWP7T $T=576120 507800 1 0 $X=575830 $Y=503590
X617 1 4 DCAP32BWP7T $T=576120 523480 1 0 $X=575830 $Y=519270
X618 1 4 DCAP32BWP7T $T=576120 531320 0 0 $X=575830 $Y=531085
X619 1 4 DCAP32BWP7T $T=576120 554840 1 0 $X=575830 $Y=550630
X620 1 4 DCAP32BWP7T $T=576120 594040 0 0 $X=575830 $Y=593805
X621 1 4 DCAP32BWP7T $T=590680 547000 1 0 $X=590390 $Y=542790
X622 1 4 DCAP32BWP7T $T=591800 570520 0 0 $X=591510 $Y=570285
X623 1 4 DCAP32BWP7T $T=618120 547000 1 0 $X=617830 $Y=542790
X624 1 4 DCAP32BWP7T $T=618120 562680 1 0 $X=617830 $Y=558470
X625 1 4 DCAP32BWP7T $T=623160 570520 0 0 $X=622870 $Y=570285
X626 1 4 DCAP32BWP7T $T=623160 578360 0 0 $X=622870 $Y=578125
X627 1 4 DCAP32BWP7T $T=640520 578360 1 0 $X=640230 $Y=574150
X628 1 4 DCAP32BWP7T $T=660120 531320 0 0 $X=659830 $Y=531085
X629 1 4 DCAP32BWP7T $T=660120 578360 0 0 $X=659830 $Y=578125
X630 1 4 DCAP32BWP7T $T=664040 492120 1 0 $X=663750 $Y=487910
X631 1 4 DCAP32BWP7T $T=664600 523480 1 0 $X=664310 $Y=519270
X632 1 4 DCAP32BWP7T $T=668520 562680 1 0 $X=668230 $Y=558470
X633 1 4 DCAP32BWP7T $T=674680 515640 1 0 $X=674390 $Y=511430
X634 1 4 DCAP32BWP7T $T=702120 507800 0 0 $X=701830 $Y=507565
X635 1 4 DCAP32BWP7T $T=702120 539160 1 0 $X=701830 $Y=534950
X636 1 4 DCAP32BWP7T $T=705480 492120 0 0 $X=705190 $Y=491885
X637 1 4 DCAP32BWP7T $T=714440 570520 0 0 $X=714150 $Y=570285
X638 1 4 DCAP32BWP7T $T=715560 515640 1 0 $X=715270 $Y=511430
X639 1 4 DCAP32BWP7T $T=717240 539160 0 0 $X=716950 $Y=538925
X640 1 4 DCAP32BWP7T $T=718360 492120 1 0 $X=718070 $Y=487910
X641 1 4 DCAP32BWP7T $T=720040 594040 0 0 $X=719750 $Y=593805
X642 1 4 DCAP32BWP7T $T=722840 554840 1 0 $X=722550 $Y=550630
X643 1 4 DCAP32BWP7T $T=725080 562680 1 0 $X=724790 $Y=558470
X644 303 298 310 295 1 4 321 FA1D0BWP7T $T=515640 515640 1 0 $X=515350 $Y=511430
X645 269 305 316 323 1 4 326 FA1D0BWP7T $T=534680 499960 1 0 $X=534390 $Y=495750
X646 309 306 338 291 1 4 337 FA1D0BWP7T $T=534680 547000 1 0 $X=534390 $Y=542790
X647 296 241 318 339 1 4 340 FA1D0BWP7T $T=534680 570520 0 0 $X=534390 $Y=570285
X648 301 312 105 336 1 4 341 FA1D0BWP7T $T=535240 586200 1 0 $X=534950 $Y=581990
X649 315 336 343 345 1 4 347 FA1D0BWP7T $T=538600 554840 0 0 $X=538310 $Y=554605
X650 334 342 352 333 1 4 356 FA1D0BWP7T $T=544200 507800 0 0 $X=543910 $Y=507565
X651 106 107 109 342 1 4 355 FA1D0BWP7T $T=544760 492120 1 0 $X=544470 $Y=487910
X652 344 348 113 361 1 4 363 FA1D0BWP7T $T=548120 586200 1 0 $X=547830 $Y=581990
X653 319 353 354 364 1 4 368 FA1D0BWP7T $T=550920 562680 1 0 $X=550630 $Y=558470
X654 356 349 369 373 1 4 374 FA1D0BWP7T $T=557080 515640 0 0 $X=556790 $Y=515405
X655 350 365 370 372 1 4 375 FA1D0BWP7T $T=557640 492120 1 0 $X=557350 $Y=487910
X656 114 355 372 369 1 4 376 FA1D0BWP7T $T=557640 499960 0 0 $X=557350 $Y=499725
X657 378 117 364 359 1 4 357 FA1D0BWP7T $T=570520 562680 1 180 $X=557350 $Y=562445
X658 314 322 283 366 1 4 379 FA1D0BWP7T $T=557640 578360 1 0 $X=557350 $Y=574150
X659 116 366 363 119 1 4 380 FA1D0BWP7T $T=557640 594040 1 0 $X=557350 $Y=589830
X660 127 397 375 384 1 4 381 FA1D0BWP7T $T=589560 499960 1 180 $X=576390 $Y=499725
X661 361 341 399 401 1 4 130 FA1D0BWP7T $T=577240 586200 0 0 $X=576950 $Y=585965
X662 347 385 401 404 1 4 131 FA1D0BWP7T $T=579480 554840 0 0 $X=579190 $Y=554605
X663 351 390 409 378 1 4 413 FA1D0BWP7T $T=586760 578360 0 0 $X=586470 $Y=578125
X664 391 132 381 418 1 4 417 FA1D0BWP7T $T=589000 507800 0 0 $X=588710 $Y=507565
X665 129 406 135 397 1 4 137 FA1D0BWP7T $T=589560 499960 1 0 $X=589270 $Y=495750
X666 367 408 420 399 1 4 140 FA1D0BWP7T $T=592360 594040 1 0 $X=592070 $Y=589830
X667 379 138 431 434 1 4 423 FA1D0BWP7T $T=599640 578360 0 0 $X=599350 $Y=578125
X668 434 359 380 159 1 4 443 FA1D0BWP7T $T=619800 594040 1 0 $X=619510 $Y=589830
X669 44 4 1 253 INVD1BWP7T $T=494920 507800 0 0 $X=494630 $Y=507565
X670 324 4 1 104 INVD1BWP7T $T=536360 554840 1 180 $X=534390 $Y=554605
X671 383 4 1 244 INVD1BWP7T $T=578360 515640 1 180 $X=576390 $Y=515405
X672 414 4 1 259 INVD1BWP7T $T=612520 562680 0 180 $X=610550 $Y=558470
X673 411 4 1 101 INVD1BWP7T $T=623160 570520 1 180 $X=621190 $Y=570285
X674 155 4 1 143 INVD1BWP7T $T=623720 507800 0 180 $X=621750 $Y=503590
X675 450 4 1 68 INVD1BWP7T $T=654520 562680 0 180 $X=652550 $Y=558470
X676 171 4 1 212 CKBD0BWP7T $T=738520 554840 1 180 $X=735990 $Y=554605
X783 7 4 11 13 1 ND2D1BWP7T $T=450680 562680 0 0 $X=450390 $Y=562445
X784 30 4 39 29 1 ND2D1BWP7T $T=461320 531320 0 0 $X=461030 $Y=531085
X785 258 4 260 63 1 ND2D1BWP7T $T=480360 539160 0 0 $X=480070 $Y=538925
X786 54 4 94 62 1 ND2D1BWP7T $T=521800 570520 1 0 $X=521510 $Y=566310
X787 98 4 102 82 1 ND2D1BWP7T $T=526280 586200 0 0 $X=525990 $Y=585965
X788 324 4 415 414 1 ND2D1BWP7T $T=596840 554840 0 0 $X=596550 $Y=554605
X789 154 4 421 112 1 ND2D1BWP7T $T=621480 492120 0 0 $X=621190 $Y=491885
X790 362 4 400 285 1 ND2D1BWP7T $T=623720 547000 0 0 $X=623430 $Y=546765
X791 398 4 435 383 1 ND2D1BWP7T $T=625960 531320 0 0 $X=625670 $Y=531085
X792 258 4 405 271 1 ND2D1BWP7T $T=628760 547000 0 0 $X=628470 $Y=546765
X793 360 4 410 63 1 ND2D1BWP7T $T=636600 594040 1 0 $X=636310 $Y=589830
X794 134 4 441 450 1 ND2D1BWP7T $T=638280 562680 1 0 $X=637990 $Y=558470
X795 307 4 438 411 1 ND2D1BWP7T $T=644440 547000 0 180 $X=641910 $Y=542790
X796 187 4 454 190 1 ND2D1BWP7T $T=666840 523480 0 0 $X=666550 $Y=523245
X797 187 4 175 192 1 ND2D1BWP7T $T=673560 523480 0 0 $X=673270 $Y=523245
X798 187 4 197 196 1 ND2D1BWP7T $T=679160 578360 0 0 $X=678870 $Y=578125
X799 194 4 500 198 1 ND2D1BWP7T $T=690920 578360 1 180 $X=688390 $Y=578125
X800 194 4 195 199 1 ND2D1BWP7T $T=688680 594040 0 0 $X=688390 $Y=593805
X801 194 4 490 200 1 ND2D1BWP7T $T=689800 539160 1 0 $X=689510 $Y=534950
X802 194 4 499 203 1 ND2D1BWP7T $T=691480 547000 0 0 $X=691190 $Y=546765
X827 247 4 1 263 INVD0BWP7T $T=484840 523480 1 0 $X=484550 $Y=519270
X828 277 4 1 279 INVD0BWP7T $T=497160 507800 0 0 $X=496870 $Y=507565
X829 270 4 1 278 INVD0BWP7T $T=501640 499960 1 180 $X=499670 $Y=499725
X830 257 4 1 284 INVD0BWP7T $T=507240 523480 1 180 $X=505270 $Y=523245
X831 234 4 1 286 INVD0BWP7T $T=505560 562680 0 0 $X=505270 $Y=562445
X832 82 4 1 81 INVD0BWP7T $T=511720 578360 0 180 $X=509750 $Y=574150
X833 292 4 1 302 INVD0BWP7T $T=521800 547000 1 180 $X=519830 $Y=546765
X834 93 4 1 96 INVD0BWP7T $T=522360 523480 0 0 $X=522070 $Y=523245
X835 308 4 1 315 INVD0BWP7T $T=525720 499960 0 0 $X=525430 $Y=499725
X836 323 4 1 310 INVD0BWP7T $T=535240 507800 0 0 $X=534950 $Y=507565
X837 326 4 1 331 INVD0BWP7T $T=536920 507800 0 0 $X=536630 $Y=507565
X838 333 4 1 329 INVD0BWP7T $T=540280 507800 1 180 $X=538310 $Y=507565
X839 95 4 1 334 INVD0BWP7T $T=539160 484280 0 0 $X=538870 $Y=484045
X840 339 4 1 338 INVD0BWP7T $T=555960 547000 1 180 $X=553990 $Y=546765
X841 337 4 1 377 INVD0BWP7T $T=568840 547000 0 0 $X=568550 $Y=546765
X842 387 4 1 391 INVD0BWP7T $T=578360 515640 1 0 $X=578070 $Y=511430
X843 41 239 44 26 4 1 OAI21D0BWP7T $T=476440 523480 1 0 $X=476150 $Y=519270
X844 288 293 289 40 4 1 OAI21D0BWP7T $T=511720 499960 0 0 $X=511430 $Y=499725
X845 290 309 282 308 4 1 OAI21D0BWP7T $T=518440 539160 0 0 $X=518150 $Y=538925
X846 92 303 83 95 4 1 OAI21D0BWP7T $T=521240 484280 0 0 $X=520950 $Y=484045
X847 325 327 321 40 4 1 OAI21D0BWP7T $T=537480 523480 0 0 $X=537190 $Y=523245
X848 396 430 374 40 4 1 OAI21D0BWP7T $T=612520 539160 1 180 $X=609430 $Y=538925
X849 448 451 168 461 4 1 OAI21D0BWP7T $T=639960 594040 1 0 $X=639670 $Y=589830
X850 448 446 454 460 4 1 OAI21D0BWP7T $T=647800 539160 1 0 $X=647510 $Y=534950
X851 174 449 175 462 4 1 OAI21D0BWP7T $T=649480 507800 0 0 $X=649190 $Y=507565
X852 175 447 176 463 4 1 OAI21D0BWP7T $T=649480 515640 0 0 $X=649190 $Y=515405
X853 448 445 175 465 4 1 OAI21D0BWP7T $T=651720 523480 0 0 $X=651430 $Y=523245
X854 454 453 176 468 4 1 OAI21D0BWP7T $T=660680 539160 1 0 $X=660390 $Y=534950
X855 181 452 454 466 4 1 OAI21D0BWP7T $T=663480 578360 0 180 $X=660390 $Y=574150
X856 174 476 454 472 4 1 OAI21D0BWP7T $T=668520 562680 0 180 $X=665430 $Y=558470
X857 184 480 454 474 4 1 OAI21D0BWP7T $T=671880 578360 0 180 $X=668790 $Y=574150
X858 191 482 454 478 4 1 OAI21D0BWP7T $T=672440 531320 0 180 $X=669350 $Y=527110
X859 448 479 195 481 4 1 OAI21D0BWP7T $T=679720 586200 1 180 $X=676630 $Y=585965
X860 191 485 175 484 4 1 OAI21D0BWP7T $T=681400 515640 1 180 $X=678310 $Y=515405
X861 448 488 490 493 4 1 OAI21D0BWP7T $T=681960 531320 0 0 $X=681670 $Y=531085
X862 448 486 197 489 4 1 OAI21D0BWP7T $T=687000 586200 1 180 $X=683910 $Y=585965
X863 448 496 499 495 4 1 OAI21D0BWP7T $T=686440 554840 0 0 $X=686150 $Y=554605
X864 490 504 176 498 4 1 OAI21D0BWP7T $T=692040 515640 1 180 $X=688950 $Y=515405
X865 448 492 500 501 4 1 OAI21D0BWP7T $T=689240 562680 1 0 $X=688950 $Y=558470
X866 175 487 181 469 4 1 OAI21D0BWP7T $T=693720 507800 1 180 $X=690630 $Y=507565
X867 197 510 176 506 4 1 OAI21D0BWP7T $T=694840 586200 1 180 $X=691750 $Y=585965
X868 174 512 490 509 4 1 OAI21D0BWP7T $T=696520 523480 1 180 $X=693430 $Y=523245
X869 499 511 176 513 4 1 OAI21D0BWP7T $T=693720 554840 1 0 $X=693430 $Y=550630
X870 500 514 176 508 4 1 OAI21D0BWP7T $T=696520 562680 1 180 $X=693430 $Y=562445
X871 174 518 500 517 4 1 OAI21D0BWP7T $T=705480 570520 1 180 $X=702390 $Y=570285
X872 191 522 490 520 4 1 OAI21D0BWP7T $T=712200 523480 1 180 $X=709110 $Y=523245
X873 174 524 499 521 4 1 OAI21D0BWP7T $T=714440 554840 1 180 $X=711350 $Y=554605
X874 184 523 490 527 4 1 OAI21D0BWP7T $T=713880 515640 0 0 $X=713590 $Y=515405
X875 191 530 500 528 4 1 OAI21D0BWP7T $T=717240 578360 1 0 $X=716950 $Y=574150
X876 184 540 500 537 4 1 OAI21D0BWP7T $T=725080 562680 0 180 $X=721990 $Y=558470
X877 184 546 499 533 4 1 OAI21D0BWP7T $T=728440 531320 1 180 $X=725350 $Y=531085
X878 191 544 499 535 4 1 OAI21D0BWP7T $T=730120 554840 1 180 $X=727030 $Y=554605
X879 499 549 181 554 4 1 OAI21D0BWP7T $T=729000 515640 0 0 $X=728710 $Y=515405
X880 205 551 213 214 4 1 OAI21D0BWP7T $T=735720 484280 0 0 $X=735430 $Y=484045
X881 490 552 181 526 4 1 OAI21D0BWP7T $T=738520 515640 0 180 $X=735430 $Y=511430
X882 500 553 181 543 4 1 OAI21D0BWP7T $T=738520 570520 1 180 $X=735430 $Y=570285
X922 43 4 54 55 1 34 ND3D0BWP7T $T=472520 586200 1 0 $X=472230 $Y=581990
X923 69 4 258 285 1 257 ND3D0BWP7T $T=504440 531320 1 0 $X=504150 $Y=527110
X924 282 4 258 307 1 308 ND3D0BWP7T $T=519560 523480 0 0 $X=519270 $Y=523245
X925 153 4 411 63 1 407 ND3D0BWP7T $T=621480 562680 1 180 $X=618390 $Y=562445
X926 170 4 145 112 1 428 ND3D0BWP7T $T=636040 492120 0 180 $X=632950 $Y=487910
X927 4 1 DCAP16BWP7T $T=450120 492120 0 0 $X=449830 $Y=491885
X928 4 1 DCAP16BWP7T $T=450120 507800 1 0 $X=449830 $Y=503590
X929 4 1 DCAP16BWP7T $T=450120 578360 1 0 $X=449830 $Y=574150
X930 4 1 DCAP16BWP7T $T=465240 578360 1 0 $X=464950 $Y=574150
X931 4 1 DCAP16BWP7T $T=472520 562680 1 0 $X=472230 $Y=558470
X932 4 1 DCAP16BWP7T $T=473080 570520 0 0 $X=472790 $Y=570285
X933 4 1 DCAP16BWP7T $T=480920 515640 0 0 $X=480630 $Y=515405
X934 4 1 DCAP16BWP7T $T=492120 499960 1 0 $X=491830 $Y=495750
X935 4 1 DCAP16BWP7T $T=492120 523480 0 0 $X=491830 $Y=523245
X936 4 1 DCAP16BWP7T $T=492120 531320 1 0 $X=491830 $Y=527110
X937 4 1 DCAP16BWP7T $T=492120 539160 0 0 $X=491830 $Y=538925
X938 4 1 DCAP16BWP7T $T=492120 578360 1 0 $X=491830 $Y=574150
X939 4 1 DCAP16BWP7T $T=494920 539160 1 0 $X=494630 $Y=534950
X940 4 1 DCAP16BWP7T $T=498840 507800 0 0 $X=498550 $Y=507565
X941 4 1 DCAP16BWP7T $T=501080 578360 0 0 $X=500790 $Y=578125
X942 4 1 DCAP16BWP7T $T=515640 492120 1 0 $X=515350 $Y=487910
X943 4 1 DCAP16BWP7T $T=521800 547000 1 0 $X=521510 $Y=542790
X944 4 1 DCAP16BWP7T $T=521800 547000 0 0 $X=521510 $Y=546765
X945 4 1 DCAP16BWP7T $T=523480 554840 1 0 $X=523190 $Y=550630
X946 4 1 DCAP16BWP7T $T=524040 570520 0 0 $X=523750 $Y=570285
X947 4 1 DCAP16BWP7T $T=534120 492120 1 0 $X=533830 $Y=487910
X948 4 1 DCAP16BWP7T $T=534120 562680 1 0 $X=533830 $Y=558470
X949 4 1 DCAP16BWP7T $T=534120 570520 1 0 $X=533830 $Y=566310
X950 4 1 DCAP16BWP7T $T=563800 562680 1 0 $X=563510 $Y=558470
X951 4 1 DCAP16BWP7T $T=576120 531320 1 0 $X=575830 $Y=527110
X952 4 1 DCAP16BWP7T $T=576120 539160 0 0 $X=575830 $Y=538925
X953 4 1 DCAP16BWP7T $T=576120 547000 1 0 $X=575830 $Y=542790
X954 4 1 DCAP16BWP7T $T=576120 562680 0 0 $X=575830 $Y=562445
X955 4 1 DCAP16BWP7T $T=576120 578360 0 0 $X=575830 $Y=578125
X956 4 1 DCAP16BWP7T $T=576120 594040 1 0 $X=575830 $Y=589830
X957 4 1 DCAP16BWP7T $T=581720 547000 0 0 $X=581430 $Y=546765
X958 4 1 DCAP16BWP7T $T=605240 539160 1 0 $X=604950 $Y=534950
X959 4 1 DCAP16BWP7T $T=618120 484280 0 0 $X=617830 $Y=484045
X960 4 1 DCAP16BWP7T $T=625960 499960 1 0 $X=625670 $Y=495750
X961 4 1 DCAP16BWP7T $T=628200 531320 0 0 $X=627910 $Y=531085
X962 4 1 DCAP16BWP7T $T=640520 562680 1 0 $X=640230 $Y=558470
X963 4 1 DCAP16BWP7T $T=641640 547000 0 0 $X=641350 $Y=546765
X964 4 1 DCAP16BWP7T $T=647240 586200 0 0 $X=646950 $Y=585965
X965 4 1 DCAP16BWP7T $T=648360 515640 1 0 $X=648070 $Y=511430
X966 4 1 DCAP16BWP7T $T=660120 554840 0 0 $X=659830 $Y=554605
X967 4 1 DCAP16BWP7T $T=680840 539160 1 0 $X=680550 $Y=534950
X968 4 1 DCAP16BWP7T $T=689240 554840 0 0 $X=688950 $Y=554605
X969 4 1 DCAP16BWP7T $T=689800 523480 1 0 $X=689510 $Y=519270
X970 4 1 DCAP16BWP7T $T=690360 570520 0 0 $X=690070 $Y=570285
X971 4 1 DCAP16BWP7T $T=690920 578360 0 0 $X=690630 $Y=578125
X972 4 1 DCAP16BWP7T $T=690920 594040 0 0 $X=690630 $Y=593805
X973 4 1 DCAP16BWP7T $T=692040 539160 1 0 $X=691750 $Y=534950
X974 4 1 DCAP16BWP7T $T=692040 562680 1 0 $X=691750 $Y=558470
X975 4 1 DCAP16BWP7T $T=702120 484280 0 0 $X=701830 $Y=484045
X976 4 1 DCAP16BWP7T $T=702120 499960 1 0 $X=701830 $Y=495750
X977 4 1 DCAP16BWP7T $T=702120 554840 0 0 $X=701830 $Y=554605
X978 4 1 DCAP16BWP7T $T=702120 586200 1 0 $X=701830 $Y=581990
X979 4 1 DCAP16BWP7T $T=712200 523480 0 0 $X=711910 $Y=523245
X980 4 1 DCAP16BWP7T $T=713320 594040 1 0 $X=713030 $Y=589830
X981 4 1 DCAP16BWP7T $T=714440 554840 0 0 $X=714150 $Y=554605
X982 4 1 DCAP16BWP7T $T=714440 562680 0 0 $X=714150 $Y=562445
X983 4 1 DCAP16BWP7T $T=722280 531320 1 0 $X=721990 $Y=527110
X984 4 1 DCAP16BWP7T $T=725640 586200 1 0 $X=725350 $Y=581990
X985 4 1 DCAP16BWP7T $T=727320 507800 0 0 $X=727030 $Y=507565
X986 4 1 DCAP16BWP7T $T=727320 570520 1 0 $X=727030 $Y=566310
X987 4 1 DCAP16BWP7T $T=729560 547000 1 0 $X=729270 $Y=542790
X1016 65 4 67 263 269 1 NR3D1BWP7T $T=482040 492120 0 0 $X=481750 $Y=491885
X1017 87 4 67 279 281 1 NR3D1BWP7T $T=521240 499960 0 0 $X=520950 $Y=499725
X1018 281 287 4 1 289 298 MAOI222D1BWP7T $T=508360 507800 0 0 $X=508070 $Y=507565
X1019 321 331 4 1 329 349 MAOI222D1BWP7T $T=547560 523480 1 0 $X=547270 $Y=519270
X1020 377 345 4 1 340 382 MAOI222D1BWP7T $T=577240 547000 0 0 $X=576950 $Y=546765
X1021 374 376 4 1 384 387 MAOI222D1BWP7T $T=589000 515640 1 180 $X=584230 $Y=515405
X1022 31 26 4 23 236 1 AOI21D1BWP7T $T=461880 562680 0 180 $X=458230 $Y=558470
X1023 289 288 4 293 274 1 AOI21D1BWP7T $T=508360 499960 0 0 $X=508070 $Y=499725
X1024 46 47 1 4 INVD2BWP7T $T=466360 531320 1 180 $X=463830 $Y=531085
X1025 26 37 1 4 INVD2BWP7T $T=499960 492120 1 0 $X=499670 $Y=487910
X1026 285 71 1 4 INVD2BWP7T $T=507800 515640 0 180 $X=505270 $Y=511430
X1027 63 48 1 4 INVD2BWP7T $T=507800 547000 0 0 $X=507510 $Y=546765
X1028 307 249 1 4 INVD2BWP7T $T=518440 562680 1 180 $X=515910 $Y=562445
X1029 258 74 1 4 INVD2BWP7T $T=519560 547000 1 0 $X=519270 $Y=542790
X1030 398 240 1 4 INVD2BWP7T $T=596840 554840 1 180 $X=594310 $Y=554605
X1083 28 230 4 1 5 DFQD0BWP7T $T=461320 531320 1 180 $X=450390 $Y=531085
X1084 28 20 4 1 228 DFQD0BWP7T $T=461320 547000 0 180 $X=450390 $Y=542790
X1085 28 21 4 1 6 DFQD0BWP7T $T=461320 554840 1 180 $X=450390 $Y=554605
X1086 28 246 4 1 35 DFQD0BWP7T $T=472520 586200 0 180 $X=461590 $Y=581990
X1087 28 248 4 1 235 DFQD0BWP7T $T=473080 570520 1 180 $X=462150 $Y=570285
X1088 28 51 4 1 45 DFQD0BWP7T $T=474760 554840 1 180 $X=463830 $Y=554605
X1089 28 53 4 1 46 DFQD0BWP7T $T=475320 594040 1 180 $X=464390 $Y=593805
X1090 28 242 4 1 238 DFQD0BWP7T $T=477000 547000 0 180 $X=466070 $Y=542790
X1091 28 256 4 1 13 DFQD0BWP7T $T=485400 570520 0 180 $X=474470 $Y=566310
X1092 28 261 4 1 58 DFQD0BWP7T $T=486520 554840 1 180 $X=475590 $Y=554605
X1093 28 266 4 1 59 DFQD0BWP7T $T=486520 594040 1 180 $X=475590 $Y=593805
X1094 28 77 4 1 70 DFQD0BWP7T $T=503320 484280 1 180 $X=492390 $Y=484045
X1095 28 274 4 1 247 DFQD0BWP7T $T=492680 531320 0 0 $X=492390 $Y=531085
X1096 28 275 4 1 282 DFQD0BWP7T $T=492680 547000 0 0 $X=492390 $Y=546765
X1097 28 280 4 1 69 DFQD0BWP7T $T=503320 562680 0 180 $X=492390 $Y=558470
X1098 28 276 4 1 277 DFQD0BWP7T $T=494360 523480 1 0 $X=494070 $Y=519270
X1099 28 251 4 1 234 DFQD0BWP7T $T=507800 570520 1 180 $X=496870 $Y=570285
X1100 28 273 4 1 272 DFQD0BWP7T $T=511160 586200 1 180 $X=500230 $Y=585965
X1101 28 300 4 1 98 DFQD0BWP7T $T=515080 594040 1 0 $X=514790 $Y=589830
X1102 28 294 4 1 83 DFQD0BWP7T $T=516200 531320 0 0 $X=515910 $Y=531085
X1103 28 335 4 1 89 DFQD0BWP7T $T=545320 594040 1 180 $X=534390 $Y=593805
X1104 28 332 4 1 317 DFQD0BWP7T $T=536360 531320 1 0 $X=536070 $Y=527110
X1105 28 346 4 1 90 DFQD0BWP7T $T=554280 570520 0 180 $X=543350 $Y=566310
X1106 28 118 4 1 362 DFQD0BWP7T $T=570520 531320 0 180 $X=559590 $Y=527110
X1107 28 371 4 1 358 DFQD0BWP7T $T=570520 539160 1 180 $X=559590 $Y=538925
X1108 28 386 4 1 398 DFQD0BWP7T $T=576680 539160 1 0 $X=576390 $Y=534950
X1109 28 388 4 1 389 DFQD0BWP7T $T=577240 523480 0 0 $X=576950 $Y=523245
X1110 28 403 4 1 411 DFQD0BWP7T $T=588440 539160 0 0 $X=588150 $Y=538925
X1111 128 412 4 1 425 DFQD0BWP7T $T=596280 523480 1 0 $X=595990 $Y=519270
X1112 128 442 4 1 437 DFQD0BWP7T $T=634360 523480 1 180 $X=623430 $Y=523245
X1113 128 444 4 1 439 DFQD0BWP7T $T=636040 515640 0 180 $X=625110 $Y=511430
X1114 128 447 4 1 456 DFQD0BWP7T $T=637160 523480 0 0 $X=636870 $Y=523245
X1115 128 165 4 1 173 DFQD0BWP7T $T=637720 499960 1 0 $X=637430 $Y=495750
X1116 128 449 4 1 457 DFQD0BWP7T $T=637720 515640 1 0 $X=637430 $Y=511430
X1117 167 452 4 1 459 DFQD0BWP7T $T=639400 562680 0 0 $X=639110 $Y=562445
X1118 128 453 4 1 458 DFQD0BWP7T $T=642200 554840 1 0 $X=641910 $Y=550630
X1119 167 455 4 1 464 DFQD0BWP7T $T=643880 578360 0 0 $X=643590 $Y=578125
X1120 128 183 4 1 483 DFQD0BWP7T $T=662360 499960 1 0 $X=662070 $Y=495750
X1121 128 480 4 1 473 DFQD0BWP7T $T=675800 562680 1 180 $X=664870 $Y=562445
X1122 128 476 4 1 471 DFQD0BWP7T $T=677480 547000 1 180 $X=666550 $Y=546765
X1123 128 482 4 1 475 DFQD0BWP7T $T=680840 539160 0 180 $X=669910 $Y=534950
X1124 128 487 4 1 467 DFQD0BWP7T $T=685880 499960 0 180 $X=674950 $Y=495750
X1125 128 485 4 1 470 DFQD0BWP7T $T=686440 507800 1 180 $X=675510 $Y=507565
X1126 128 504 4 1 494 DFQD0BWP7T $T=696520 499960 1 180 $X=685590 $Y=499725
X1127 167 510 4 1 491 DFQD0BWP7T $T=713320 594040 0 180 $X=702390 $Y=589830
X1128 128 518 4 1 503 DFQD0BWP7T $T=713880 578360 1 180 $X=702950 $Y=578125
X1129 128 522 4 1 507 DFQD0BWP7T $T=714440 499960 1 180 $X=703510 $Y=499725
X1130 128 514 4 1 505 DFQD0BWP7T $T=714440 562680 1 180 $X=703510 $Y=562445
X1131 128 523 4 1 516 DFQD0BWP7T $T=715560 515640 0 180 $X=704630 $Y=511430
X1132 128 512 4 1 502 DFQD0BWP7T $T=715560 531320 0 180 $X=704630 $Y=527110
X1133 128 511 4 1 497 DFQD0BWP7T $T=715560 554840 0 180 $X=704630 $Y=550630
X1134 128 524 4 1 515 DFQD0BWP7T $T=717240 539160 1 180 $X=706310 $Y=538925
X1135 128 530 4 1 525 DFQD0BWP7T $T=725640 586200 0 180 $X=714710 $Y=581990
X1136 128 534 4 1 542 DFQD0BWP7T $T=717800 499960 1 0 $X=717510 $Y=495750
X1137 128 544 4 1 531 DFQD0BWP7T $T=729560 547000 0 180 $X=718630 $Y=542790
X1138 167 550 4 1 541 DFQD0BWP7T $T=734600 594040 0 180 $X=723670 $Y=589830
X1139 128 552 4 1 529 DFQD0BWP7T $T=738520 507800 0 180 $X=727590 $Y=503590
X1140 128 549 4 1 538 DFQD0BWP7T $T=738520 523480 0 180 $X=727590 $Y=519270
X1141 128 539 4 1 547 DFQD0BWP7T $T=738520 539160 0 180 $X=727590 $Y=534950
X1142 128 546 4 1 536 DFQD0BWP7T $T=738520 547000 1 180 $X=727590 $Y=546765
X1143 128 540 4 1 532 DFQD0BWP7T $T=738520 562680 1 180 $X=727590 $Y=562445
X1144 128 553 4 1 548 DFQD0BWP7T $T=738520 578360 1 180 $X=727590 $Y=578125
X1145 44 4 1 37 33 237 NR3D0BWP7T $T=464120 507800 0 180 $X=461030 $Y=503590
X1146 44 4 1 37 33 264 NR3D0BWP7T $T=480920 499960 1 0 $X=480630 $Y=495750
X1147 286 4 1 74 48 296 NR3D0BWP7T $T=506120 562680 1 0 $X=505830 $Y=558470
X1148 270 267 264 52 4 1 AOI21D0BWP7T $T=484280 499960 1 180 $X=481190 $Y=499725
X1149 97 304 263 269 4 1 AOI21D0BWP7T $T=525720 499960 0 180 $X=522630 $Y=495750
X1150 325 332 321 327 4 1 AOI21D0BWP7T $T=539160 515640 1 180 $X=536070 $Y=515405
X1151 396 426 374 430 4 1 AOI21D0BWP7T $T=612520 523480 1 180 $X=609430 $Y=523245
X1152 62 60 4 1 56 AN2D1BWP7T $T=478120 578360 0 180 $X=475030 $Y=574150
X1153 271 60 4 1 261 AN2D1BWP7T $T=484280 547000 0 180 $X=481190 $Y=542790
X1154 90 60 4 1 84 AN2D1BWP7T $T=516200 578360 1 180 $X=513110 $Y=578125
X1155 89 60 4 1 91 AN2D1BWP7T $T=517880 586200 0 0 $X=517590 $Y=585965
X1156 360 60 4 1 335 AN2D1BWP7T $T=567720 547000 1 180 $X=564630 $Y=546765
X1157 362 60 4 1 346 AN2D1BWP7T $T=590680 547000 0 180 $X=587590 $Y=542790
X1158 373 40 4 1 388 AN2D1BWP7T $T=603000 539160 0 0 $X=602710 $Y=538925
X1159 360 285 4 1 353 AN2D1BWP7T $T=621480 554840 0 180 $X=618390 $Y=550630
X1160 418 40 4 1 442 AN2D1BWP7T $T=660680 554840 1 0 $X=660390 $Y=550630
X1161 345 340 337 1 4 313 XOR3D0BWP7T $T=552040 539160 1 180 $X=542230 $Y=538925
X1162 284 302 299 1 4 252 XNR3D0BWP7T $T=523480 554840 0 180 $X=513670 $Y=550630
X1163 253 270 4 66 1 262 267 OAI22D1BWP7T $T=486520 507800 0 180 $X=482310 $Y=503590
X1164 24 277 4 280 255 1 IOA21D0BWP7T $T=496040 515640 0 0 $X=495750 $Y=515405
X1165 34 4 40 43 1 49 42 OAI211D0BWP7T $T=461880 578360 1 0 $X=461590 $Y=574150
X1166 257 4 40 69 1 254 255 OAI211D0BWP7T $T=480920 531320 1 180 $X=477270 $Y=531085
X1167 389 40 404 24 4 1 133 AO22D0BWP7T $T=591800 547000 0 0 $X=591510 $Y=546765
X1168 284 299 302 306 4 1 MAOI222D2BWP7T $T=512280 523480 0 0 $X=511990 $Y=523245
X1169 28 22 4 1 8 DFQD1BWP7T $T=461320 570520 1 180 $X=450390 $Y=570285
X1170 28 233 4 1 9 DFQD1BWP7T $T=461320 586200 0 180 $X=450390 $Y=581990
X1171 28 262 4 1 44 DFQD1BWP7T $T=485960 531320 0 180 $X=475030 $Y=527110
X1172 28 64 4 1 57 DFQD1BWP7T $T=486520 492120 0 180 $X=475590 $Y=487910
X1173 28 311 4 1 115 DFQD1BWP7T $T=548120 547000 1 0 $X=547830 $Y=542790
X1174 28 330 4 1 324 DFQD1BWP7T $T=549240 531320 1 0 $X=548950 $Y=527110
X1175 128 402 4 1 134 DFQD1BWP7T $T=587880 531320 1 0 $X=587590 $Y=527110
X1176 128 426 4 1 136 DFQD1BWP7T $T=610280 531320 1 180 $X=599350 $Y=531085
X1177 128 440 4 1 151 DFQD1BWP7T $T=629320 539160 0 180 $X=618390 $Y=534950
X1178 128 445 4 1 383 DFQD1BWP7T $T=641640 539160 0 180 $X=630710 $Y=534950
X1179 128 446 4 1 271 DFQD1BWP7T $T=641640 547000 1 180 $X=630710 $Y=546765
X1180 167 451 4 1 414 DFQD1BWP7T $T=647240 586200 1 180 $X=636310 $Y=585965
X1181 167 479 4 1 182 DFQD1BWP7T $T=673000 586200 1 180 $X=662070 $Y=585965
X1182 128 486 4 1 450 DFQD1BWP7T $T=684760 578360 0 180 $X=673830 $Y=574150
X1183 128 488 4 1 307 DFQD1BWP7T $T=686440 523480 1 180 $X=675510 $Y=523245
X1184 128 201 4 1 477 DFQD1BWP7T $T=695400 492120 0 180 $X=684470 $Y=487910
X1185 128 206 4 1 519 DFQD1BWP7T $T=718360 492120 0 180 $X=707430 $Y=487910
X1186 128 551 4 1 545 DFQD1BWP7T $T=738520 492120 1 180 $X=727590 $Y=491885
X1187 24 234 4 1 19 18 17 MOAI22D0BWP7T $T=459080 594040 1 180 $X=454870 $Y=593805
X1188 24 282 4 1 79 266 19 MOAI22D0BWP7T $T=510040 594040 0 180 $X=505830 $Y=589830
X1189 24 317 4 1 313 311 19 MOAI22D0BWP7T $T=528520 523480 1 180 $X=524310 $Y=523245
X1190 24 169 4 1 19 440 427 MOAI22D0BWP7T $T=643320 531320 1 180 $X=639110 $Y=531085
X1191 10 14 231 25 36 4 1 XNR4D0BWP7T $T=450680 499960 1 0 $X=450390 $Y=495750
X1192 407 410 416 419 423 4 1 XNR4D0BWP7T $T=592920 562680 0 0 $X=592630 $Y=562445
X1193 416 415 427 395 433 4 1 XNR4D0BWP7T $T=599080 554840 1 0 $X=598790 $Y=550630
X1194 148 428 422 421 417 4 1 XNR4D0BWP7T $T=612520 507800 0 180 $X=599350 $Y=503590
X1195 38 27 229 15 5 4 1 XOR4D0BWP7T $T=463560 507800 1 180 $X=450390 $Y=507565
X1196 405 400 395 124 357 4 1 XOR4D0BWP7T $T=591800 570520 1 180 $X=578630 $Y=570285
X1197 435 438 419 441 163 4 1 XOR4D0BWP7T $T=621480 562680 0 0 $X=621190 $Y=562445
X1198 368 413 433 443 151 4 1 XOR4D0BWP7T $T=627640 578360 1 0 $X=627350 $Y=574150
X1199 154 4 1 392 CKND1BWP7T $T=621480 492120 1 180 $X=619510 $Y=491885
X1200 170 4 1 142 CKND1BWP7T $T=643880 492120 1 180 $X=641910 $Y=491885
X1201 235 32 4 1 BUFFD1P5BWP7T $T=459080 578360 1 0 $X=458790 $Y=574150
X1202 172 55 4 1 BUFFD1P5BWP7T $T=648920 492120 0 180 $X=645830 $Y=487910
X1203 477 188 4 1 BUFFD1P5BWP7T $T=670200 484280 1 180 $X=667110 $Y=484045
X1204 519 204 4 1 BUFFD1P5BWP7T $T=705480 492120 1 180 $X=702390 $Y=491885
X1205 545 211 4 1 BUFFD1P5BWP7T $T=727320 484280 1 180 $X=724230 $Y=484045
X1206 249 1 23 248 4 NR2D0BWP7T $T=472520 562680 0 180 $X=469990 $Y=558470
X1207 326 329 1 331 4 333 325 AOI22D1BWP7T $T=536360 515640 1 0 $X=536070 $Y=511430
X1208 228 4 1 12 CKBD1BWP7T $T=450680 547000 0 0 $X=450390 $Y=546765
X1209 238 4 1 29 CKBD1BWP7T $T=462440 523480 0 180 $X=459910 $Y=519270
X1210 272 4 1 54 CKBD1BWP7T $T=483720 570520 0 0 $X=483430 $Y=570285
X1211 358 4 1 360 CKBD1BWP7T $T=557640 539160 0 0 $X=557350 $Y=538925
X1212 425 4 1 152 CKBD1BWP7T $T=620920 547000 1 180 $X=618390 $Y=546765
X1213 437 4 1 145 CKBD1BWP7T $T=639400 562680 1 180 $X=636870 $Y=562445
X1214 439 4 1 169 CKBD1BWP7T $T=651720 531320 1 180 $X=649190 $Y=531085
X1215 287 281 1 4 281 288 287 MAOI22D0BWP7T $T=511720 499960 0 180 $X=507510 $Y=495750
X1216 464 171 1 4 171 455 454 MAOI22D0BWP7T $T=649480 570520 1 180 $X=645270 $Y=570285
X1217 542 171 1 4 212 534 490 MAOI22D0BWP7T $T=727320 507800 1 180 $X=723110 $Y=507565
X1218 547 171 1 4 212 539 499 MAOI22D0BWP7T $T=727320 523480 1 180 $X=723110 $Y=523245
X1219 541 171 1 4 212 550 500 MAOI22D0BWP7T $T=734600 594040 1 0 $X=734310 $Y=589830
X1220 429 145 428 1 4 150 OA21D0BWP7T $T=609160 492120 1 0 $X=608870 $Y=487910
X1221 153 436 407 1 4 431 OA21D0BWP7T $T=621480 578360 1 0 $X=621190 $Y=574150
X1222 458 460 271 178 448 1 4 AOI22D0BWP7T $T=647800 547000 1 0 $X=647510 $Y=542790
X1223 180 461 414 178 448 1 4 AOI22D0BWP7T $T=654520 594040 0 180 $X=650870 $Y=589830
X1224 181 469 178 467 173 1 4 AOI22D0BWP7T $T=664040 492120 0 180 $X=660390 $Y=487910
X1225 174 462 178 457 470 1 4 AOI22D0BWP7T $T=660680 507800 0 0 $X=660390 $Y=507565
X1226 181 466 178 459 464 1 4 AOI22D0BWP7T $T=660680 570520 1 0 $X=660390 $Y=566310
X1227 176 463 178 456 457 1 4 AOI22D0BWP7T $T=664600 523480 0 180 $X=660950 $Y=519270
X1228 176 468 178 458 471 1 4 AOI22D0BWP7T $T=661240 539160 0 0 $X=660950 $Y=538925
X1229 456 465 383 178 448 1 4 AOI22D0BWP7T $T=665160 531320 0 180 $X=661510 $Y=527110
X1230 174 472 178 471 475 1 4 AOI22D0BWP7T $T=664040 554840 1 0 $X=663750 $Y=550630
X1231 184 474 178 473 459 1 4 AOI22D0BWP7T $T=667960 578360 0 180 $X=664310 $Y=574150
X1232 184 185 178 483 467 1 4 AOI22D0BWP7T $T=665160 499960 0 0 $X=664870 $Y=499725
X1233 191 478 178 475 473 1 4 AOI22D0BWP7T $T=670200 539160 0 180 $X=666550 $Y=534950
X1234 193 481 182 178 448 1 4 AOI22D0BWP7T $T=671880 594040 0 180 $X=668230 $Y=589830
X1235 191 484 178 470 483 1 4 AOI22D0BWP7T $T=671320 515640 1 0 $X=671030 $Y=511430
X1236 491 489 450 178 448 1 4 AOI22D0BWP7T $T=684200 586200 1 180 $X=680550 $Y=585965
X1237 497 495 285 178 448 1 4 AOI22D0BWP7T $T=687000 539160 1 180 $X=683350 $Y=538925
X1238 494 493 307 178 448 1 4 AOI22D0BWP7T $T=686440 523480 1 0 $X=686150 $Y=519270
X1239 176 498 178 494 502 1 4 AOI22D0BWP7T $T=686440 531320 0 0 $X=686150 $Y=531085
X1240 505 501 63 178 448 1 4 AOI22D0BWP7T $T=690360 570520 1 180 $X=686710 $Y=570285
X1241 176 508 178 505 503 1 4 AOI22D0BWP7T $T=694280 578360 0 180 $X=690630 $Y=574150
X1242 176 506 178 491 202 1 4 AOI22D0BWP7T $T=690920 594040 1 0 $X=690630 $Y=589830
X1243 174 509 178 502 507 1 4 AOI22D0BWP7T $T=696520 531320 1 180 $X=692870 $Y=531085
X1244 176 513 178 497 515 1 4 AOI22D0BWP7T $T=693160 539160 0 0 $X=692870 $Y=538925
X1245 191 520 178 507 516 1 4 AOI22D0BWP7T $T=706040 515640 1 180 $X=702390 $Y=515405
X1246 174 521 178 515 531 1 4 AOI22D0BWP7T $T=705480 547000 1 0 $X=705190 $Y=542790
X1247 174 517 178 503 525 1 4 AOI22D0BWP7T $T=711080 570520 0 0 $X=710790 $Y=570285
X1248 209 208 204 207 205 1 4 AOI22D0BWP7T $T=718360 484280 1 180 $X=714710 $Y=484045
X1249 181 526 178 529 542 1 4 AOI22D0BWP7T $T=715560 507800 1 0 $X=715270 $Y=503590
X1250 191 528 178 525 532 1 4 AOI22D0BWP7T $T=716120 570520 1 0 $X=715830 $Y=566310
X1251 184 527 178 516 529 1 4 AOI22D0BWP7T $T=717800 515640 0 0 $X=717510 $Y=515405
X1252 184 533 178 536 538 1 4 AOI22D0BWP7T $T=718920 531320 1 0 $X=718630 $Y=527110
X1253 191 535 178 531 536 1 4 AOI22D0BWP7T $T=719480 554840 1 0 $X=719190 $Y=550630
X1254 184 537 178 532 548 1 4 AOI22D0BWP7T $T=723960 570520 1 0 $X=723670 $Y=566310
X1255 181 543 178 548 541 1 4 AOI22D0BWP7T $T=724520 578360 1 0 $X=724230 $Y=574150
X1256 181 554 178 538 547 1 4 AOI22D0BWP7T $T=735160 531320 1 0 $X=734870 $Y=527110
X1257 4 1 ICV_41 $T=468040 507800 1 0 $X=467750 $Y=503590
X1258 4 1 ICV_41 $T=468040 515640 1 0 $X=467750 $Y=511430
X1259 4 1 ICV_41 $T=492120 515640 1 0 $X=491830 $Y=511430
X1260 4 1 ICV_41 $T=503320 484280 0 0 $X=503030 $Y=484045
X1261 4 1 ICV_41 $T=518440 492120 0 0 $X=518150 $Y=491885
X1262 4 1 ICV_41 $T=576120 499960 1 0 $X=575830 $Y=495750
X1263 4 1 ICV_41 $T=589000 492120 1 0 $X=588710 $Y=487910
X1264 4 1 ICV_41 $T=589000 515640 0 0 $X=588710 $Y=515405
X1265 4 1 ICV_41 $T=618120 492120 1 0 $X=617830 $Y=487910
X1266 4 1 ICV_41 $T=643880 507800 1 0 $X=643590 $Y=503590
X1267 4 1 ICV_41 $T=644440 523480 1 0 $X=644150 $Y=519270
X1268 4 1 ICV_41 $T=685880 499960 1 0 $X=685590 $Y=495750
X1269 4 1 ICV_41 $T=702120 507800 1 0 $X=701830 $Y=503590
X1270 4 1 ICV_41 $T=702120 570520 1 0 $X=701830 $Y=566310
X1271 4 1 ICV_41 $T=702120 594040 0 0 $X=701830 $Y=593805
X1272 4 1 ICV_41 $T=713880 578360 0 0 $X=713590 $Y=578125
X1273 4 1 ICV_41 $T=728440 531320 0 0 $X=728150 $Y=531085
X1274 4 1 ICV_37 $T=477000 539160 0 0 $X=476710 $Y=538925
X1275 4 1 ICV_37 $T=501080 531320 1 0 $X=500790 $Y=527110
X1276 4 1 ICV_37 $T=501080 539160 0 0 $X=500790 $Y=538925
X1277 4 1 ICV_37 $T=510040 578360 0 0 $X=509750 $Y=578125
X1278 4 1 ICV_37 $T=517320 499960 0 0 $X=517030 $Y=499725
X1279 4 1 ICV_37 $T=534120 523480 0 0 $X=533830 $Y=523245
X1280 4 1 ICV_37 $T=540280 507800 0 0 $X=539990 $Y=507565
X1281 4 1 ICV_37 $T=576120 554840 0 0 $X=575830 $Y=554605
X1282 4 1 ICV_37 $T=585080 539160 0 0 $X=584790 $Y=538925
X1283 4 1 ICV_37 $T=613640 484280 0 0 $X=613350 $Y=484045
X1284 4 1 ICV_37 $T=618120 570520 0 0 $X=617830 $Y=570285
X1285 4 1 ICV_37 $T=632680 594040 1 0 $X=632390 $Y=589830
X1286 4 1 ICV_37 $T=644440 547000 1 0 $X=644150 $Y=542790
X1287 4 1 ICV_37 $T=649480 562680 1 0 $X=649190 $Y=558470
X1288 4 1 ICV_37 $T=655640 547000 1 0 $X=655350 $Y=542790
X1289 4 1 ICV_37 $T=660120 515640 1 0 $X=659830 $Y=511430
X1290 4 1 ICV_37 $T=673000 586200 0 0 $X=672710 $Y=585965
X1291 4 1 ICV_37 $T=702120 547000 1 0 $X=701830 $Y=542790
X1292 4 1 ICV_37 $T=711080 484280 0 0 $X=710790 $Y=484045
X1293 4 1 ICV_37 $T=715560 531320 1 0 $X=715270 $Y=527110
X1294 4 1 ICV_37 $T=720040 507800 0 0 $X=719750 $Y=507565
X1295 4 1 ICV_37 $T=723400 554840 0 0 $X=723110 $Y=554605
X1296 4 1 ICV_37 $T=724520 547000 0 0 $X=724230 $Y=546765
X1297 4 1 ICV_37 $T=725640 515640 0 0 $X=725350 $Y=515405
X1298 4 1 ICV_37 $T=732360 570520 0 0 $X=732070 $Y=570285
X1299 4 1 ICV_43 $T=450120 523480 1 0 $X=449830 $Y=519270
X1300 4 1 ICV_43 $T=461320 547000 1 0 $X=461030 $Y=542790
X1301 4 1 ICV_43 $T=461320 554840 0 0 $X=461030 $Y=554605
X1302 4 1 ICV_43 $T=492120 507800 0 0 $X=491830 $Y=507565
X1303 4 1 ICV_43 $T=503320 562680 1 0 $X=503030 $Y=558470
X1304 4 1 ICV_43 $T=507240 562680 0 0 $X=506950 $Y=562445
X1305 4 1 ICV_43 $T=519000 570520 1 0 $X=518710 $Y=566310
X1306 4 1 ICV_43 $T=534120 484280 0 0 $X=533830 $Y=484045
X1307 4 1 ICV_43 $T=576120 570520 0 0 $X=575830 $Y=570285
X1308 4 1 ICV_43 $T=585080 531320 1 0 $X=584790 $Y=527110
X1309 4 1 ICV_43 $T=585080 547000 1 0 $X=584790 $Y=542790
X1310 4 1 ICV_43 $T=618120 578360 0 0 $X=617830 $Y=578125
X1311 4 1 ICV_43 $T=620920 547000 0 0 $X=620630 $Y=546765
X1312 4 1 ICV_43 $T=624840 578360 1 0 $X=624550 $Y=574150
X1313 4 1 ICV_43 $T=634360 523480 0 0 $X=634070 $Y=523245
X1314 4 1 ICV_43 $T=634360 562680 0 0 $X=634070 $Y=562445
X1315 4 1 ICV_43 $T=634920 499960 1 0 $X=634630 $Y=495750
X1316 4 1 ICV_43 $T=639400 554840 1 0 $X=639110 $Y=550630
X1317 4 1 ICV_43 $T=641080 578360 0 0 $X=640790 $Y=578125
X1318 4 1 ICV_43 $T=673000 507800 0 0 $X=672710 $Y=507565
X1319 4 1 ICV_43 $T=681960 492120 1 0 $X=681670 $Y=487910
X1320 4 1 ICV_43 $T=685880 578360 0 0 $X=685590 $Y=578125
X1321 4 1 ICV_43 $T=686440 562680 1 0 $X=686150 $Y=558470
X1322 4 1 ICV_43 $T=702120 515640 1 0 $X=701830 $Y=511430
X1323 4 1 ICV_43 $T=702120 531320 1 0 $X=701830 $Y=527110
X1324 4 1 ICV_43 $T=702120 554840 1 0 $X=701830 $Y=550630
X1325 4 1 ICV_55 $T=468040 492120 1 0 $X=467750 $Y=487910
X1326 4 1 ICV_55 $T=492120 492120 1 0 $X=491830 $Y=487910
X1327 4 1 ICV_55 $T=507800 570520 0 0 $X=507510 $Y=570285
X1328 4 1 ICV_55 $T=525160 531320 1 0 $X=524870 $Y=527110
X1329 4 1 ICV_55 $T=543080 562680 1 0 $X=542790 $Y=558470
X1330 4 1 ICV_55 $T=567160 515640 1 0 $X=566870 $Y=511430
X1331 4 1 ICV_55 $T=567160 523480 0 0 $X=566870 $Y=523245
X1332 4 1 ICV_55 $T=585080 562680 0 0 $X=584790 $Y=562445
X1333 4 1 ICV_55 $T=603000 562680 1 0 $X=602710 $Y=558470
X1334 4 1 ICV_55 $T=618120 531320 0 0 $X=617830 $Y=531085
X1335 4 1 ICV_55 $T=627080 484280 0 0 $X=626790 $Y=484045
X1336 4 1 ICV_55 $T=678600 554840 0 0 $X=678310 $Y=554605
X1337 4 1 ICV_55 $T=681400 515640 0 0 $X=681110 $Y=515405
X1338 4 1 ICV_55 $T=706040 515640 0 0 $X=705750 $Y=515405
X1339 4 1 ICV_55 $T=720040 523480 1 0 $X=719750 $Y=519270
X1340 4 1 ICV_55 $T=720040 539160 1 0 $X=719750 $Y=534950
X1341 4 1 ICV_55 $T=735160 539160 0 0 $X=734870 $Y=538925
X1342 4 1 ICV_54 $T=459080 594040 0 0 $X=458790 $Y=593805
X1343 4 1 ICV_54 $T=485400 515640 1 0 $X=485110 $Y=511430
X1344 4 1 ICV_54 $T=485400 562680 1 0 $X=485110 $Y=558470
X1345 4 1 ICV_54 $T=485400 570520 1 0 $X=485110 $Y=566310
X1346 4 1 ICV_54 $T=500520 594040 1 0 $X=500230 $Y=589830
X1347 4 1 ICV_54 $T=504440 578360 1 0 $X=504150 $Y=574150
X1348 4 1 ICV_54 $T=513960 547000 1 0 $X=513670 $Y=542790
X1349 4 1 ICV_54 $T=527400 562680 0 0 $X=527110 $Y=562445
X1350 4 1 ICV_54 $T=552040 539160 0 0 $X=551750 $Y=538925
X1351 4 1 ICV_54 $T=552040 562680 0 0 $X=551750 $Y=562445
X1352 4 1 ICV_54 $T=552040 578360 1 0 $X=551750 $Y=574150
X1353 4 1 ICV_54 $T=552040 594040 1 0 $X=551750 $Y=589830
X1354 4 1 ICV_54 $T=569400 554840 0 0 $X=569110 $Y=554605
X1355 4 1 ICV_54 $T=594040 507800 1 0 $X=593750 $Y=503590
X1356 4 1 ICV_54 $T=594040 531320 0 0 $X=593750 $Y=531085
X1357 4 1 ICV_54 $T=618120 523480 0 0 $X=617830 $Y=523245
X1358 4 1 ICV_54 $T=660120 562680 1 0 $X=659830 $Y=558470
X1359 4 1 ICV_54 $T=688120 562680 0 0 $X=687830 $Y=562445
X1360 4 1 ICV_54 $T=695400 492120 1 0 $X=695110 $Y=487910
X1361 4 1 ICV_54 $T=702120 492120 1 0 $X=701830 $Y=487910
X1362 4 1 ICV_54 $T=737400 499960 1 0 $X=737110 $Y=495750
X1363 4 1 ICV_38 $T=486520 492120 1 0 $X=486230 $Y=487910
X1364 4 1 ICV_38 $T=486520 492120 0 0 $X=486230 $Y=491885
X1365 4 1 ICV_38 $T=486520 554840 0 0 $X=486230 $Y=554605
X1366 4 1 ICV_38 $T=486520 586200 1 0 $X=486230 $Y=581990
X1367 4 1 ICV_38 $T=486520 594040 0 0 $X=486230 $Y=593805
X1368 4 1 ICV_38 $T=528520 507800 1 0 $X=528230 $Y=503590
X1369 4 1 ICV_38 $T=528520 515640 1 0 $X=528230 $Y=511430
X1370 4 1 ICV_38 $T=528520 523480 0 0 $X=528230 $Y=523245
X1371 4 1 ICV_38 $T=528520 562680 1 0 $X=528230 $Y=558470
X1372 4 1 ICV_38 $T=528520 586200 1 0 $X=528230 $Y=581990
X1373 4 1 ICV_38 $T=528520 586200 0 0 $X=528230 $Y=585965
X1374 4 1 ICV_38 $T=570520 492120 1 0 $X=570230 $Y=487910
X1375 4 1 ICV_38 $T=570520 499960 0 0 $X=570230 $Y=499725
X1376 4 1 ICV_38 $T=570520 531320 1 0 $X=570230 $Y=527110
X1377 4 1 ICV_38 $T=570520 539160 0 0 $X=570230 $Y=538925
X1378 4 1 ICV_38 $T=570520 562680 0 0 $X=570230 $Y=562445
X1379 4 1 ICV_38 $T=570520 578360 1 0 $X=570230 $Y=574150
X1380 4 1 ICV_38 $T=570520 594040 1 0 $X=570230 $Y=589830
X1381 4 1 ICV_38 $T=612520 492120 1 0 $X=612230 $Y=487910
X1382 4 1 ICV_38 $T=612520 507800 1 0 $X=612230 $Y=503590
X1383 4 1 ICV_38 $T=612520 523480 0 0 $X=612230 $Y=523245
X1384 4 1 ICV_38 $T=612520 539160 0 0 $X=612230 $Y=538925
X1385 4 1 ICV_38 $T=612520 562680 1 0 $X=612230 $Y=558470
X1386 4 1 ICV_38 $T=612520 562680 0 0 $X=612230 $Y=562445
X1387 4 1 ICV_38 $T=612520 594040 1 0 $X=612230 $Y=589830
X1388 4 1 ICV_38 $T=612520 594040 0 0 $X=612230 $Y=593805
X1389 4 1 ICV_38 $T=654520 523480 0 0 $X=654230 $Y=523245
X1390 4 1 ICV_38 $T=654520 562680 1 0 $X=654230 $Y=558470
X1391 4 1 ICV_38 $T=654520 594040 1 0 $X=654230 $Y=589830
X1392 4 1 ICV_38 $T=696520 499960 0 0 $X=696230 $Y=499725
X1393 4 1 ICV_38 $T=696520 523480 0 0 $X=696230 $Y=523245
X1394 4 1 ICV_38 $T=696520 539160 0 0 $X=696230 $Y=538925
X1395 4 1 ICV_38 $T=696520 554840 1 0 $X=696230 $Y=550630
X1396 4 1 ICV_38 $T=738520 484280 0 0 $X=738230 $Y=484045
X1397 4 1 ICV_38 $T=738520 492120 0 0 $X=738230 $Y=491885
X1398 4 1 ICV_38 $T=738520 507800 1 0 $X=738230 $Y=503590
X1399 4 1 ICV_38 $T=738520 515640 1 0 $X=738230 $Y=511430
X1400 4 1 ICV_38 $T=738520 523480 1 0 $X=738230 $Y=519270
X1401 4 1 ICV_38 $T=738520 531320 1 0 $X=738230 $Y=527110
X1402 4 1 ICV_38 $T=738520 539160 1 0 $X=738230 $Y=534950
X1403 4 1 ICV_38 $T=738520 547000 1 0 $X=738230 $Y=542790
X1404 4 1 ICV_38 $T=738520 547000 0 0 $X=738230 $Y=546765
X1405 4 1 ICV_38 $T=738520 554840 0 0 $X=738230 $Y=554605
X1406 4 1 ICV_38 $T=738520 562680 0 0 $X=738230 $Y=562445
X1407 4 1 ICV_38 $T=738520 570520 0 0 $X=738230 $Y=570285
X1408 4 1 ICV_38 $T=738520 578360 0 0 $X=738230 $Y=578125
X1409 4 1 ICV_38 $T=738520 594040 1 0 $X=738230 $Y=589830
X1410 4 1 ICV_45 $T=450120 539160 0 0 $X=449830 $Y=538925
X1411 4 1 ICV_45 $T=463560 507800 0 0 $X=463270 $Y=507565
X1412 4 1 ICV_45 $T=492120 570520 1 0 $X=491830 $Y=566310
X1413 4 1 ICV_45 $T=492120 586200 1 0 $X=491830 $Y=581990
X1414 4 1 ICV_45 $T=499400 515640 0 0 $X=499110 $Y=515405
X1415 4 1 ICV_45 $T=501640 507800 1 0 $X=501350 $Y=503590
X1416 4 1 ICV_45 $T=540280 515640 1 0 $X=539990 $Y=511430
X1417 4 1 ICV_45 $T=540280 523480 0 0 $X=539990 $Y=523245
X1418 4 1 ICV_45 $T=545320 594040 0 0 $X=545030 $Y=593805
X1419 4 1 ICV_45 $T=576120 562680 1 0 $X=575830 $Y=558470
X1420 4 1 ICV_45 $T=589560 499960 0 0 $X=589270 $Y=499725
X1421 4 1 ICV_45 $T=620920 515640 0 0 $X=620630 $Y=515405
X1422 4 1 ICV_45 $T=660120 570520 0 0 $X=659830 $Y=570285
X1423 4 1 ICV_45 $T=660120 594040 0 0 $X=659830 $Y=593805
X1424 4 1 ICV_45 $T=670200 484280 0 0 $X=669910 $Y=484045
X1425 4 1 ICV_45 $T=672440 531320 1 0 $X=672150 $Y=527110
X1426 4 1 ICV_45 $T=714440 499960 0 0 $X=714150 $Y=499725
X1427 239 4 1 31 BUFFD3BWP7T $T=463560 523480 1 0 $X=463270 $Y=519270
X1428 237 4 1 50 BUFFD3BWP7T $T=464120 507800 1 0 $X=463830 $Y=503590
X1429 243 4 1 52 BUFFD3BWP7T $T=468040 499960 1 0 $X=467750 $Y=495750
X1430 210 4 1 200 BUFFD3BWP7T $T=720040 594040 1 180 $X=715830 $Y=593805
X1431 304 4 1 289 BUFFD1BWP7T $T=517320 499960 1 180 $X=514790 $Y=499725
X1432 187 4 1 194 BUFFD1BWP7T $T=678600 554840 1 180 $X=676070 $Y=554605
X1433 317 320 4 1 350 352 IAO21D0BWP7T $T=553720 499960 0 0 $X=553430 $Y=499725
X1434 115 328 4 1 367 343 IAO21D0BWP7T $T=564360 547000 1 180 $X=560710 $Y=546765
X1435 389 123 4 1 120 365 IAO21D0BWP7T $T=580040 492120 0 180 $X=576390 $Y=487910
X1436 136 424 4 1 139 406 IAO21D0BWP7T $T=606920 492120 0 180 $X=603270 $Y=487910
X1437 146 147 4 1 144 408 IAO21D0BWP7T $T=612520 594040 1 180 $X=608870 $Y=593805
X1438 112 111 317 1 4 350 AN3D1BWP7T $T=557080 499960 0 180 $X=553430 $Y=495750
X1439 112 126 389 1 4 120 AN3D1BWP7T $T=589000 492120 0 180 $X=585350 $Y=487910
X1440 63 324 115 1 4 367 AN3D1BWP7T $T=610280 562680 1 180 $X=606630 $Y=562445
X1441 63 134 146 1 4 144 AN3D1BWP7T $T=612520 594040 0 180 $X=608870 $Y=589830
X1442 112 155 136 1 4 139 AN3D1BWP7T $T=638280 484280 1 180 $X=634630 $Y=484045
X1443 28 61 41 4 1 DFQD2BWP7T $T=480920 515640 1 180 $X=469430 $Y=515405
X1444 28 268 258 4 1 DFQD2BWP7T $T=504440 539160 0 0 $X=504150 $Y=538925
X1445 128 492 63 4 1 DFQD2BWP7T $T=688120 562680 1 180 $X=676630 $Y=562445
X1446 128 496 285 4 1 DFQD2BWP7T $T=689800 547000 1 180 $X=678310 $Y=546765
X1447 141 156 4 1 BUFFD2BWP7T $T=622600 499960 1 0 $X=622310 $Y=495750
X1448 161 162 164 4 1 ND2D2BWP7T $T=630440 507800 1 0 $X=630150 $Y=503590
X1449 177 179 164 4 1 ND2D2BWP7T $T=650040 499960 1 0 $X=649750 $Y=495750
X1450 158 448 166 4 1 ND2D1P5BWP7T $T=639960 507800 1 0 $X=639670 $Y=503590
X1451 24 247 4 19 251 252 1 MOAI22D1BWP7T $T=469160 531320 0 0 $X=468870 $Y=531085
X1452 24 83 4 291 275 19 1 MOAI22D1BWP7T $T=513400 523480 0 180 $X=508630 $Y=519270
X1453 232 1 16 231 4 230 229 AOI211D1BWP7T $T=456280 523480 0 180 $X=452630 $Y=519270
X1454 19 1 281 76 4 276 279 AOI211D1BWP7T $T=501640 507800 0 180 $X=497990 $Y=503590
X1455 432 1 19 422 4 444 149 AOI211D1BWP7T $T=620920 507800 0 0 $X=620630 $Y=507565
X1456 72 28 4 1 INVD10BWP7T $T=492680 578360 0 0 $X=492390 $Y=578125
X1457 86 72 4 1 INVD10BWP7T $T=515640 570520 0 0 $X=515350 $Y=570285
X1479 164 186 189 4 1 INR2XD2BWP7T $T=663480 515640 1 0 $X=663190 $Y=511430
X1480 41 278 75 33 270 1 4 73 OA32D0BWP7T $T=499960 499960 1 180 $X=494070 $Y=499725
X1481 236 40 4 1 BUFFD6BWP7T $T=493800 594040 1 0 $X=493510 $Y=589830
X1482 85 4 270 80 78 37 1 OAI31D2BWP7T $T=515640 492120 0 180 $X=508630 $Y=487910
X1483 164 4 160 158 1 ND2D3BWP7T $T=635480 492120 1 180 $X=630150 $Y=491885
X1484 382 4 1 385 CKND0BWP7T $T=576680 515640 1 0 $X=576390 $Y=511430
.ENDS
***************************************
.SUBCKT ICV_48 1 2
** N=2 EP=2 IP=4 FDC=34
*.SEEDPROM
X0 1 2 ICV_40 $T=17920 0 0 0 $X=17630 $Y=-235
X1 2 1 DCAP32BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_53 2 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175
** N=626 EP=173 IP=5057 FDC=13734
*.SEEDPROM
M0 6 64 221 6 N L=1.8e-07 W=5e-07 $X=476500 $Y=655780 $D=0
M1 623 223 6 6 N L=1.8e-07 W=5e-07 $X=477285 $Y=655415 $D=0
M2 226 64 623 6 N L=1.8e-07 W=5e-07 $X=477905 $Y=655780 $D=0
M3 223 221 226 6 N L=1.8e-07 W=5e-07 $X=478705 $Y=655780 $D=0
M4 6 214 223 6 N L=1.8e-07 W=1e-06 $X=479465 $Y=655415 $D=0
M5 6 226 231 6 N L=1.8e-07 W=5e-07 $X=480995 $Y=655800 $D=0
M6 624 235 6 6 N L=1.8e-07 W=5e-07 $X=481795 $Y=655415 $D=0
M7 239 231 624 6 N L=1.8e-07 W=5e-07 $X=482225 $Y=655415 $D=0
M8 235 226 239 6 N L=1.8e-07 W=5e-07 $X=483085 $Y=655820 $D=0
M9 6 213 235 6 N L=1.8e-07 W=1e-06 $X=483845 $Y=655415 $D=0
M10 243 239 6 6 N L=1.8e-07 W=1e-06 $X=484595 $Y=655415 $D=0
M11 5 64 221 5 P L=1.8e-07 W=6.85e-07 $X=476500 $Y=653280 $D=16
M12 625 223 5 5 P L=1.8e-07 W=6.85e-07 $X=477285 $Y=653650 $D=16
M13 226 221 625 5 P L=1.8e-07 W=6.85e-07 $X=477865 $Y=653650 $D=16
M14 223 64 226 5 P L=1.8e-07 W=6.85e-07 $X=478665 $Y=653650 $D=16
M15 5 214 223 5 P L=1.8e-07 W=1.37e-06 $X=479425 $Y=653185 $D=16
M16 5 226 231 5 P L=1.8e-07 W=6.85e-07 $X=480995 $Y=653260 $D=16
M17 626 235 5 5 P L=1.8e-07 W=6.85e-07 $X=481795 $Y=653630 $D=16
M18 239 226 626 5 P L=1.8e-07 W=6.85e-07 $X=482305 $Y=653630 $D=16
M19 235 231 239 5 P L=1.8e-07 W=6.85e-07 $X=483045 $Y=653630 $D=16
M20 5 213 235 5 P L=1.8e-07 W=1.37e-06 $X=483825 $Y=653185 $D=16
M21 243 239 5 5 P L=1.8e-07 W=1.37e-06 $X=484595 $Y=653185 $D=16
X34 4 5 6 6 2 174 175 175 174 622 174 6 PDDW0208CDG $T=900240 610000 0 90 $X=780240 $Y=609400
X228 5 6 DCAPBWP7T $T=450120 648920 1 0 $X=449830 $Y=644710
X229 5 6 DCAPBWP7T $T=454600 688120 0 0 $X=454310 $Y=687885
X230 5 6 DCAPBWP7T $T=456840 625400 1 0 $X=456550 $Y=621190
X231 5 6 DCAPBWP7T $T=478120 625400 0 0 $X=477830 $Y=625165
X232 5 6 DCAPBWP7T $T=480920 609720 1 0 $X=480630 $Y=605510
X233 5 6 DCAPBWP7T $T=482600 735160 1 0 $X=482310 $Y=730950
X234 5 6 DCAPBWP7T $T=489320 601880 0 0 $X=489030 $Y=601645
X235 5 6 DCAPBWP7T $T=489320 633240 1 0 $X=489030 $Y=629030
X236 5 6 DCAPBWP7T $T=489320 695960 0 0 $X=489030 $Y=695725
X237 5 6 DCAPBWP7T $T=489320 727320 1 0 $X=489030 $Y=723110
X238 5 6 DCAPBWP7T $T=498840 672440 1 0 $X=498550 $Y=668230
X239 5 6 DCAPBWP7T $T=498840 672440 0 0 $X=498550 $Y=672205
X240 5 6 DCAPBWP7T $T=513960 641080 0 0 $X=513670 $Y=640845
X241 5 6 DCAPBWP7T $T=534120 641080 0 0 $X=533830 $Y=640845
X242 5 6 DCAPBWP7T $T=534120 735160 0 0 $X=533830 $Y=734925
X243 5 6 DCAPBWP7T $T=544200 633240 0 0 $X=543910 $Y=633005
X244 5 6 DCAPBWP7T $T=544760 601880 1 0 $X=544470 $Y=597670
X245 5 6 DCAPBWP7T $T=573320 719480 0 0 $X=573030 $Y=719245
X246 5 6 DCAPBWP7T $T=573320 735160 0 0 $X=573030 $Y=734925
X247 5 6 DCAPBWP7T $T=576120 711640 1 0 $X=575830 $Y=707430
X248 5 6 DCAPBWP7T $T=578920 601880 1 0 $X=578630 $Y=597670
X249 5 6 DCAPBWP7T $T=589560 656760 1 0 $X=589270 $Y=652550
X250 5 6 DCAPBWP7T $T=591800 617560 0 0 $X=591510 $Y=617325
X251 5 6 DCAPBWP7T $T=597960 625400 0 0 $X=597670 $Y=625165
X252 5 6 DCAPBWP7T $T=600200 617560 0 0 $X=599910 $Y=617325
X253 5 6 DCAPBWP7T $T=604120 727320 1 0 $X=603830 $Y=723110
X254 5 6 DCAPBWP7T $T=607480 711640 0 0 $X=607190 $Y=711405
X255 5 6 DCAPBWP7T $T=615320 641080 0 0 $X=615030 $Y=640845
X256 5 6 DCAPBWP7T $T=615320 703800 1 0 $X=615030 $Y=699590
X257 5 6 DCAPBWP7T $T=615320 727320 1 0 $X=615030 $Y=723110
X258 5 6 DCAPBWP7T $T=618120 601880 0 0 $X=617830 $Y=601645
X259 5 6 DCAPBWP7T $T=625400 641080 0 0 $X=625110 $Y=640845
X260 5 6 DCAPBWP7T $T=631000 735160 0 0 $X=630710 $Y=734925
X261 5 6 DCAPBWP7T $T=639400 711640 1 0 $X=639110 $Y=707430
X262 5 6 DCAPBWP7T $T=642200 641080 0 0 $X=641910 $Y=640845
X263 5 6 DCAPBWP7T $T=642760 664600 1 0 $X=642470 $Y=660390
X264 5 6 DCAPBWP7T $T=649480 719480 0 0 $X=649190 $Y=719245
X265 5 6 DCAPBWP7T $T=657320 695960 0 0 $X=657030 $Y=695725
X266 5 6 DCAPBWP7T $T=660120 680280 0 0 $X=659830 $Y=680045
X267 5 6 DCAPBWP7T $T=666840 727320 1 0 $X=666550 $Y=723110
X268 5 6 DCAPBWP7T $T=676920 680280 0 0 $X=676630 $Y=680045
X269 5 6 DCAPBWP7T $T=679720 664600 0 0 $X=679430 $Y=664365
X270 5 6 DCAPBWP7T $T=681960 703800 0 0 $X=681670 $Y=703565
X271 5 6 DCAPBWP7T $T=683080 625400 0 0 $X=682790 $Y=625165
X272 5 6 DCAPBWP7T $T=684760 727320 0 0 $X=684470 $Y=727085
X273 5 6 DCAPBWP7T $T=691480 617560 0 0 $X=691190 $Y=617325
X274 5 6 DCAPBWP7T $T=699320 609720 1 0 $X=699030 $Y=605510
X275 5 6 DCAPBWP7T $T=699320 648920 0 0 $X=699030 $Y=648685
X276 5 6 DCAPBWP7T $T=706600 617560 1 0 $X=706310 $Y=613350
X277 5 6 DCAPBWP7T $T=708840 617560 0 0 $X=708550 $Y=617325
X278 5 6 DCAPBWP7T $T=715560 648920 1 0 $X=715270 $Y=644710
X279 5 6 DCAPBWP7T $T=717800 719480 1 0 $X=717510 $Y=715270
X280 5 6 DCAPBWP7T $T=726200 680280 0 0 $X=725910 $Y=680045
X281 5 6 DCAPBWP7T $T=727320 617560 0 0 $X=727030 $Y=617325
X282 5 6 DCAPBWP7T $T=732360 719480 1 0 $X=732070 $Y=715270
X283 5 6 DCAPBWP7T $T=734040 688120 0 0 $X=733750 $Y=687885
X284 5 6 DCAPBWP7T $T=741320 625400 0 0 $X=741030 $Y=625165
X285 5 6 DCAPBWP7T $T=741320 648920 1 0 $X=741030 $Y=644710
X286 5 6 DCAPBWP7T $T=741320 695960 1 0 $X=741030 $Y=691750
X287 6 5 DCAP8BWP7T $T=450120 688120 0 0 $X=449830 $Y=687885
X288 6 5 DCAP8BWP7T $T=452920 672440 1 0 $X=452630 $Y=668230
X289 6 5 DCAP8BWP7T $T=466920 617560 1 0 $X=466630 $Y=613350
X290 6 5 DCAP8BWP7T $T=471960 648920 1 0 $X=471670 $Y=644710
X291 6 5 DCAP8BWP7T $T=484840 633240 1 0 $X=484550 $Y=629030
X292 6 5 DCAP8BWP7T $T=484840 688120 0 0 $X=484550 $Y=687885
X293 6 5 DCAP8BWP7T $T=484840 695960 0 0 $X=484550 $Y=695725
X294 6 5 DCAP8BWP7T $T=507800 601880 0 0 $X=507510 $Y=601645
X295 6 5 DCAP8BWP7T $T=510040 719480 1 0 $X=509750 $Y=715270
X296 6 5 DCAP8BWP7T $T=526840 695960 1 0 $X=526550 $Y=691750
X297 6 5 DCAP8BWP7T $T=527960 648920 1 0 $X=527670 $Y=644710
X298 6 5 DCAP8BWP7T $T=528520 672440 1 0 $X=528230 $Y=668230
X299 6 5 DCAP8BWP7T $T=528520 711640 1 0 $X=528230 $Y=707430
X300 6 5 DCAP8BWP7T $T=534120 633240 0 0 $X=533830 $Y=633005
X301 6 5 DCAP8BWP7T $T=534120 695960 0 0 $X=533830 $Y=695725
X302 6 5 DCAP8BWP7T $T=552040 601880 0 0 $X=551750 $Y=601645
X303 6 5 DCAP8BWP7T $T=552040 680280 0 0 $X=551750 $Y=680045
X304 6 5 DCAP8BWP7T $T=568840 727320 0 0 $X=568550 $Y=727085
X305 6 5 DCAP8BWP7T $T=568840 735160 0 0 $X=568550 $Y=734925
X306 6 5 DCAP8BWP7T $T=568840 743000 1 0 $X=568550 $Y=738790
X307 6 5 DCAP8BWP7T $T=569400 656760 0 0 $X=569110 $Y=656525
X308 6 5 DCAP8BWP7T $T=569960 633240 1 0 $X=569670 $Y=629030
X309 6 5 DCAP8BWP7T $T=570520 601880 0 0 $X=570230 $Y=601645
X310 6 5 DCAP8BWP7T $T=576120 695960 0 0 $X=575830 $Y=695725
X311 6 5 DCAP8BWP7T $T=576120 727320 0 0 $X=575830 $Y=727085
X312 6 5 DCAP8BWP7T $T=589560 656760 0 0 $X=589270 $Y=656525
X313 6 5 DCAP8BWP7T $T=592360 680280 0 0 $X=592070 $Y=680045
X314 6 5 DCAP8BWP7T $T=595720 617560 0 0 $X=595430 $Y=617325
X315 6 5 DCAP8BWP7T $T=601320 688120 0 0 $X=601030 $Y=687885
X316 6 5 DCAP8BWP7T $T=611400 601880 1 0 $X=611110 $Y=597670
X317 6 5 DCAP8BWP7T $T=611400 672440 0 0 $X=611110 $Y=672205
X318 6 5 DCAP8BWP7T $T=611400 727320 0 0 $X=611110 $Y=727085
X319 6 5 DCAP8BWP7T $T=612520 656760 1 0 $X=612230 $Y=652550
X320 6 5 DCAP8BWP7T $T=612520 664600 0 0 $X=612230 $Y=664365
X321 6 5 DCAP8BWP7T $T=618120 688120 0 0 $X=617830 $Y=687885
X322 6 5 DCAP8BWP7T $T=618120 719480 1 0 $X=617830 $Y=715270
X323 6 5 DCAP8BWP7T $T=620920 641080 0 0 $X=620630 $Y=640845
X324 6 5 DCAP8BWP7T $T=629320 727320 1 0 $X=629030 $Y=723110
X325 6 5 DCAP8BWP7T $T=634360 680280 0 0 $X=634070 $Y=680045
X326 6 5 DCAP8BWP7T $T=636040 641080 1 0 $X=635750 $Y=636870
X327 6 5 DCAP8BWP7T $T=641080 727320 1 0 $X=640790 $Y=723110
X328 6 5 DCAP8BWP7T $T=643320 688120 1 0 $X=643030 $Y=683910
X329 6 5 DCAP8BWP7T $T=652840 601880 1 0 $X=652550 $Y=597670
X330 6 5 DCAP8BWP7T $T=652840 648920 0 0 $X=652550 $Y=648685
X331 6 5 DCAP8BWP7T $T=652840 703800 1 0 $X=652550 $Y=699590
X332 6 5 DCAP8BWP7T $T=652840 719480 1 0 $X=652550 $Y=715270
X333 6 5 DCAP8BWP7T $T=653960 672440 1 0 $X=653670 $Y=668230
X334 6 5 DCAP8BWP7T $T=653960 680280 0 0 $X=653670 $Y=680045
X335 6 5 DCAP8BWP7T $T=654520 735160 0 0 $X=654230 $Y=734925
X336 6 5 DCAP8BWP7T $T=672440 680280 0 0 $X=672150 $Y=680045
X337 6 5 DCAP8BWP7T $T=687560 609720 0 0 $X=687270 $Y=609485
X338 6 5 DCAP8BWP7T $T=687560 664600 1 0 $X=687270 $Y=660390
X339 6 5 DCAP8BWP7T $T=694840 719480 0 0 $X=694550 $Y=719245
X340 6 5 DCAP8BWP7T $T=695400 625400 0 0 $X=695110 $Y=625165
X341 6 5 DCAP8BWP7T $T=696520 633240 0 0 $X=696230 $Y=633005
X342 6 5 DCAP8BWP7T $T=702120 617560 1 0 $X=701830 $Y=613350
X343 6 5 DCAP8BWP7T $T=702120 625400 0 0 $X=701830 $Y=625165
X344 6 5 DCAP8BWP7T $T=702120 695960 1 0 $X=701830 $Y=691750
X345 6 5 DCAP8BWP7T $T=702120 711640 1 0 $X=701830 $Y=707430
X346 6 5 DCAP8BWP7T $T=718360 625400 0 0 $X=718070 $Y=625165
X347 6 5 DCAP8BWP7T $T=729560 688120 0 0 $X=729270 $Y=687885
X348 6 5 DCAP8BWP7T $T=737400 743000 1 0 $X=737110 $Y=738790
X349 6 5 DCAP8BWP7T $T=737960 656760 1 0 $X=737670 $Y=652550
X350 6 5 DCAP8BWP7T $T=737960 719480 1 0 $X=737670 $Y=715270
X351 6 5 DCAP4BWP7T $T=470280 664600 1 0 $X=469990 $Y=660390
X352 6 5 DCAP4BWP7T $T=487080 625400 1 0 $X=486790 $Y=621190
X353 6 5 DCAP4BWP7T $T=488200 688120 1 0 $X=487910 $Y=683910
X354 6 5 DCAP4BWP7T $T=488200 703800 0 0 $X=487910 $Y=703565
X355 6 5 DCAP4BWP7T $T=488200 711640 0 0 $X=487910 $Y=711405
X356 6 5 DCAP4BWP7T $T=494920 719480 0 0 $X=494630 $Y=719245
X357 6 5 DCAP4BWP7T $T=497160 656760 1 0 $X=496870 $Y=652550
X358 6 5 DCAP4BWP7T $T=510040 719480 0 0 $X=509750 $Y=719245
X359 6 5 DCAP4BWP7T $T=523480 711640 0 0 $X=523190 $Y=711405
X360 6 5 DCAP4BWP7T $T=530200 601880 0 0 $X=529910 $Y=601645
X361 6 5 DCAP4BWP7T $T=530200 617560 0 0 $X=529910 $Y=617325
X362 6 5 DCAP4BWP7T $T=530200 656760 1 0 $X=529910 $Y=652550
X363 6 5 DCAP4BWP7T $T=530760 609720 1 0 $X=530470 $Y=605510
X364 6 5 DCAP4BWP7T $T=563240 735160 0 0 $X=562950 $Y=734925
X365 6 5 DCAP4BWP7T $T=576120 695960 1 0 $X=575830 $Y=691750
X366 6 5 DCAP4BWP7T $T=613080 735160 0 0 $X=612790 $Y=734925
X367 6 5 DCAP4BWP7T $T=614200 617560 1 0 $X=613910 $Y=613350
X368 6 5 DCAP4BWP7T $T=618120 711640 0 0 $X=617830 $Y=711405
X369 6 5 DCAP4BWP7T $T=618120 735160 0 0 $X=617830 $Y=734925
X370 6 5 DCAP4BWP7T $T=622040 656760 1 0 $X=621750 $Y=652550
X371 6 5 DCAP4BWP7T $T=656200 664600 1 0 $X=655910 $Y=660390
X372 6 5 DCAP4BWP7T $T=656760 609720 1 0 $X=656470 $Y=605510
X373 6 5 DCAP4BWP7T $T=656760 617560 1 0 $X=656470 $Y=613350
X374 6 5 DCAP4BWP7T $T=656760 633240 1 0 $X=656470 $Y=629030
X375 6 5 DCAP4BWP7T $T=660120 601880 1 0 $X=659830 $Y=597670
X376 6 5 DCAP4BWP7T $T=660120 656760 1 0 $X=659830 $Y=652550
X377 6 5 DCAP4BWP7T $T=673000 656760 1 0 $X=672710 $Y=652550
X378 6 5 DCAP4BWP7T $T=676360 601880 1 0 $X=676070 $Y=597670
X379 6 5 DCAP4BWP7T $T=676360 695960 1 0 $X=676070 $Y=691750
X380 6 5 DCAP4BWP7T $T=685880 656760 1 0 $X=685590 $Y=652550
X381 6 5 DCAP4BWP7T $T=688120 601880 0 0 $X=687830 $Y=601645
X382 6 5 DCAP4BWP7T $T=691480 633240 0 0 $X=691190 $Y=633005
X383 6 5 DCAP4BWP7T $T=697080 641080 1 0 $X=696790 $Y=636870
X384 6 5 DCAP4BWP7T $T=698200 601880 1 0 $X=697910 $Y=597670
X385 6 5 DCAP4BWP7T $T=698200 617560 1 0 $X=697910 $Y=613350
X386 6 5 DCAP4BWP7T $T=698760 625400 1 0 $X=698470 $Y=621190
X387 6 5 DCAP4BWP7T $T=698760 703800 1 0 $X=698470 $Y=699590
X388 6 5 DCAP4BWP7T $T=698760 703800 0 0 $X=698470 $Y=703565
X389 6 5 DCAP4BWP7T $T=698760 727320 0 0 $X=698470 $Y=727085
X390 6 5 DCAP4BWP7T $T=702120 688120 1 0 $X=701830 $Y=683910
X391 6 5 DCAP4BWP7T $T=711640 695960 0 0 $X=711350 $Y=695725
X392 6 5 DCAP4BWP7T $T=714440 609720 1 0 $X=714150 $Y=605510
X393 6 5 DCAP4BWP7T $T=740760 703800 0 0 $X=740470 $Y=703565
X394 6 5 ICV_40 $T=450120 625400 1 0 $X=449830 $Y=621190
X395 6 5 ICV_40 $T=477000 641080 1 0 $X=476710 $Y=636870
X396 6 5 ICV_40 $T=482600 727320 1 0 $X=482310 $Y=723110
X397 6 5 ICV_40 $T=483160 711640 1 0 $X=482870 $Y=707430
X398 6 5 ICV_40 $T=483720 664600 1 0 $X=483430 $Y=660390
X399 6 5 ICV_40 $T=492120 641080 1 0 $X=491830 $Y=636870
X400 6 5 ICV_40 $T=492120 672440 1 0 $X=491830 $Y=668230
X401 6 5 ICV_40 $T=492120 672440 0 0 $X=491830 $Y=672205
X402 6 5 ICV_40 $T=525720 664600 0 0 $X=525430 $Y=664365
X403 6 5 ICV_40 $T=548120 617560 1 0 $X=547830 $Y=613350
X404 6 5 ICV_40 $T=553720 719480 0 0 $X=553430 $Y=719245
X405 6 5 ICV_40 $T=561000 617560 0 0 $X=560710 $Y=617325
X406 6 5 ICV_40 $T=561000 703800 1 0 $X=560710 $Y=699590
X407 6 5 ICV_40 $T=567720 711640 1 0 $X=567430 $Y=707430
X408 6 5 ICV_40 $T=567720 711640 0 0 $X=567430 $Y=711405
X409 6 5 ICV_40 $T=568280 617560 1 0 $X=567990 $Y=613350
X410 6 5 ICV_40 $T=597400 727320 1 0 $X=597110 $Y=723110
X411 6 5 ICV_40 $T=598520 601880 0 0 $X=598230 $Y=601645
X412 6 5 ICV_40 $T=600760 711640 0 0 $X=600470 $Y=711405
X413 6 5 ICV_40 $T=608600 680280 1 0 $X=608310 $Y=676070
X414 6 5 ICV_40 $T=608600 727320 1 0 $X=608310 $Y=723110
X415 6 5 ICV_40 $T=609160 688120 0 0 $X=608870 $Y=687885
X416 6 5 ICV_40 $T=610280 625400 0 0 $X=609990 $Y=625165
X417 6 5 ICV_40 $T=610280 688120 1 0 $X=609990 $Y=683910
X418 6 5 ICV_40 $T=618120 727320 0 0 $X=617830 $Y=727085
X419 6 5 ICV_40 $T=620920 617560 1 0 $X=620630 $Y=613350
X420 6 5 ICV_40 $T=627080 633240 0 0 $X=626790 $Y=633005
X421 6 5 ICV_40 $T=634360 719480 1 0 $X=634070 $Y=715270
X422 6 5 ICV_40 $T=636600 672440 1 0 $X=636310 $Y=668230
X423 6 5 ICV_40 $T=639400 695960 0 0 $X=639110 $Y=695725
X424 6 5 ICV_40 $T=639960 601880 1 0 $X=639670 $Y=597670
X425 6 5 ICV_40 $T=645000 703800 0 0 $X=644710 $Y=703565
X426 6 5 ICV_40 $T=650600 695960 0 0 $X=650310 $Y=695725
X427 6 5 ICV_40 $T=651720 688120 1 0 $X=651430 $Y=683910
X428 6 5 ICV_40 $T=651720 711640 1 0 $X=651430 $Y=707430
X429 6 5 ICV_40 $T=660120 727320 1 0 $X=659830 $Y=723110
X430 6 5 ICV_40 $T=676920 609720 0 0 $X=676630 $Y=609485
X431 6 5 ICV_40 $T=681400 672440 0 0 $X=681110 $Y=672205
X432 6 5 ICV_40 $T=693160 601880 0 0 $X=692870 $Y=601645
X433 6 5 ICV_40 $T=693160 648920 1 0 $X=692870 $Y=644710
X434 6 5 ICV_40 $T=693160 735160 0 0 $X=692870 $Y=734925
X435 6 5 ICV_40 $T=702120 617560 0 0 $X=701830 $Y=617325
X436 6 5 ICV_40 $T=702120 664600 0 0 $X=701830 $Y=664365
X437 6 5 ICV_40 $T=702120 695960 0 0 $X=701830 $Y=695725
X438 6 5 ICV_40 $T=735720 664600 1 0 $X=735430 $Y=660390
X439 6 5 ICV_40 $T=736280 617560 1 0 $X=735990 $Y=613350
X440 187 5 181 10 6 NR2D1BWP7T $T=452920 609720 1 180 $X=450390 $Y=609485
X441 179 5 184 23 6 NR2D1BWP7T $T=450680 672440 1 0 $X=450390 $Y=668230
X442 14 5 185 24 6 NR2D1BWP7T $T=450680 688120 1 0 $X=450390 $Y=683910
X443 24 5 183 180 6 NR2D1BWP7T $T=452920 711640 0 180 $X=450390 $Y=707430
X444 22 5 189 28 6 NR2D1BWP7T $T=451800 648920 1 0 $X=451510 $Y=644710
X445 180 5 192 20 6 NR2D1BWP7T $T=457400 735160 0 0 $X=457110 $Y=734925
X446 20 5 195 32 6 NR2D1BWP7T $T=459640 735160 0 0 $X=459350 $Y=734925
X447 44 5 196 46 6 NR2D1BWP7T $T=461880 735160 0 0 $X=461590 $Y=734925
X448 180 5 201 46 6 NR2D1BWP7T $T=464120 735160 0 0 $X=463830 $Y=734925
X449 187 5 203 23 6 NR2D1BWP7T $T=465240 695960 0 0 $X=464950 $Y=695725
X450 14 5 202 53 6 NR2D1BWP7T $T=466360 735160 0 0 $X=466070 $Y=734925
X451 32 5 208 46 6 NR2D1BWP7T $T=472520 735160 1 180 $X=469990 $Y=734925
X452 180 5 216 53 6 NR2D1BWP7T $T=474760 735160 1 180 $X=472230 $Y=734925
X453 23 5 63 10 6 NR2D1BWP7T $T=477000 633240 1 180 $X=474470 $Y=633005
X454 187 5 220 68 6 NR2D1BWP7T $T=476440 648920 1 0 $X=476150 $Y=644710
X455 187 5 70 22 6 NR2D1BWP7T $T=480360 601880 1 180 $X=477830 $Y=601645
X456 224 5 71 10 6 NR2D1BWP7T $T=480920 641080 1 180 $X=478390 $Y=640845
X457 229 5 75 10 6 NR2D1BWP7T $T=483160 641080 1 180 $X=480630 $Y=640845
X458 22 5 211 179 6 NR2D1BWP7T $T=484840 609720 0 180 $X=482310 $Y=605510
X459 179 5 241 224 6 NR2D1BWP7T $T=486520 625400 1 180 $X=483990 $Y=625165
X460 247 5 78 10 6 NR2D1BWP7T $T=486520 641080 1 180 $X=483990 $Y=640845
X461 82 5 79 80 6 NR2D1BWP7T $T=494920 601880 1 180 $X=492390 $Y=601645
X462 68 5 253 179 6 NR2D1BWP7T $T=492680 609720 1 0 $X=492390 $Y=605510
X463 256 5 251 229 6 NR2D1BWP7T $T=494920 648920 1 180 $X=492390 $Y=648685
X464 179 5 254 247 6 NR2D1BWP7T $T=492680 656760 1 0 $X=492390 $Y=652550
X465 22 5 81 10 6 NR2D1BWP7T $T=494920 695960 1 180 $X=492390 $Y=695725
X466 14 5 252 69 6 NR2D1BWP7T $T=492680 727320 1 0 $X=492390 $Y=723110
X467 187 5 263 229 6 NR2D1BWP7T $T=494920 656760 1 0 $X=494630 $Y=652550
X468 14 5 261 92 6 NR2D1BWP7T $T=494920 727320 1 0 $X=494630 $Y=723110
X469 22 5 264 256 6 NR2D1BWP7T $T=498280 641080 0 0 $X=497990 $Y=640845
X470 22 5 267 266 6 NR2D1BWP7T $T=499400 656760 1 0 $X=499110 $Y=652550
X471 82 5 86 87 6 NR2D1BWP7T $T=500520 601880 0 0 $X=500230 $Y=601645
X472 23 5 271 273 6 NR2D1BWP7T $T=500520 641080 1 0 $X=500230 $Y=636870
X473 187 5 268 247 6 NR2D1BWP7T $T=502760 672440 0 180 $X=500230 $Y=668230
X474 28 5 265 10 6 NR2D1BWP7T $T=502760 672440 1 180 $X=500230 $Y=672205
X475 187 5 282 90 6 NR2D1BWP7T $T=505560 601880 0 0 $X=505270 $Y=601645
X476 22 5 283 273 6 NR2D1BWP7T $T=506120 648920 0 0 $X=505830 $Y=648685
X477 44 5 304 53 6 NR2D1BWP7T $T=526280 743000 0 180 $X=523750 $Y=738790
X478 266 5 328 224 6 NR2D1BWP7T $T=525720 711640 0 0 $X=525430 $Y=711405
X479 266 5 330 10 6 NR2D1BWP7T $T=526280 695960 0 0 $X=525990 $Y=695725
X480 273 5 331 10 6 NR2D1BWP7T $T=526280 711640 1 0 $X=525990 $Y=707430
X481 256 5 353 10 6 NR2D1BWP7T $T=542520 719480 0 0 $X=542230 $Y=719245
X482 23 5 355 256 6 NR2D1BWP7T $T=543080 695960 1 0 $X=542790 $Y=691750
X483 179 5 365 229 6 NR2D1BWP7T $T=548680 719480 1 0 $X=548390 $Y=715270
X484 179 5 367 10 6 NR2D1BWP7T $T=549240 727320 1 0 $X=548950 $Y=723110
X485 69 5 279 44 6 NR2D1BWP7T $T=552600 735160 0 0 $X=552310 $Y=734925
X486 28 5 295 247 6 NR2D1BWP7T $T=555960 695960 1 180 $X=553430 $Y=695725
X487 273 5 372 224 6 NR2D1BWP7T $T=555960 719480 0 180 $X=553430 $Y=715270
X488 28 5 378 229 6 NR2D1BWP7T $T=555960 695960 0 0 $X=555670 $Y=695725
X489 28 5 381 224 6 NR2D1BWP7T $T=560440 695960 1 180 $X=557910 $Y=695725
X490 256 5 390 224 6 NR2D1BWP7T $T=564360 719480 1 180 $X=561830 $Y=719245
X491 110 5 368 10 6 NR2D1BWP7T $T=576680 601880 1 0 $X=576390 $Y=597670
X492 134 5 132 131 6 NR2D1BWP7T $T=620920 617560 0 180 $X=618390 $Y=613350
X493 109 5 449 131 6 NR2D1BWP7T $T=620920 617560 1 180 $X=618390 $Y=617325
X494 134 5 395 10 6 NR2D1BWP7T $T=620920 641080 1 180 $X=618390 $Y=640845
X495 5 6 DCAP64BWP7T $T=452360 703800 0 0 $X=452070 $Y=703565
X496 5 6 DCAP64BWP7T $T=494920 609720 1 0 $X=494630 $Y=605510
X497 5 6 DCAP64BWP7T $T=580600 695960 1 0 $X=580310 $Y=691750
X498 5 6 DCAP64BWP7T $T=706040 601880 1 0 $X=705750 $Y=597670
X555 6 5 ICV_47 $T=450120 656760 0 0 $X=449830 $Y=656525
X556 6 5 ICV_47 $T=450120 664600 0 0 $X=449830 $Y=664365
X557 6 5 ICV_47 $T=450120 680280 0 0 $X=449830 $Y=680045
X558 6 5 ICV_47 $T=450120 727320 0 0 $X=449830 $Y=727085
X559 6 5 ICV_47 $T=492120 609720 0 0 $X=491830 $Y=609485
X560 6 5 ICV_47 $T=492120 625400 1 0 $X=491830 $Y=621190
X561 6 5 ICV_47 $T=492120 656760 0 0 $X=491830 $Y=656525
X562 6 5 ICV_47 $T=492120 664600 1 0 $X=491830 $Y=660390
X563 6 5 ICV_47 $T=492120 688120 1 0 $X=491830 $Y=683910
X564 6 5 ICV_47 $T=492120 703800 1 0 $X=491830 $Y=699590
X565 6 5 ICV_47 $T=492120 727320 0 0 $X=491830 $Y=727085
X566 6 5 ICV_47 $T=534120 609720 1 0 $X=533830 $Y=605510
X567 6 5 ICV_47 $T=534120 625400 1 0 $X=533830 $Y=621190
X568 6 5 ICV_47 $T=534120 648920 1 0 $X=533830 $Y=644710
X569 6 5 ICV_47 $T=534120 664600 1 0 $X=533830 $Y=660390
X570 6 5 ICV_47 $T=534120 672440 0 0 $X=533830 $Y=672205
X571 6 5 ICV_47 $T=534120 680280 1 0 $X=533830 $Y=676070
X572 6 5 ICV_47 $T=534120 688120 0 0 $X=533830 $Y=687885
X573 6 5 ICV_47 $T=534120 703800 0 0 $X=533830 $Y=703565
X574 6 5 ICV_47 $T=534120 735160 1 0 $X=533830 $Y=730950
X575 6 5 ICV_47 $T=576120 625400 1 0 $X=575830 $Y=621190
X576 6 5 ICV_47 $T=576120 648920 1 0 $X=575830 $Y=644710
X577 6 5 ICV_47 $T=576120 648920 0 0 $X=575830 $Y=648685
X578 6 5 ICV_47 $T=576120 664600 1 0 $X=575830 $Y=660390
X579 6 5 ICV_47 $T=576120 743000 1 0 $X=575830 $Y=738790
X580 6 5 ICV_47 $T=618120 625400 1 0 $X=617830 $Y=621190
X581 6 5 ICV_47 $T=618120 672440 0 0 $X=617830 $Y=672205
X582 6 5 ICV_47 $T=618120 735160 1 0 $X=617830 $Y=730950
X583 6 5 ICV_47 $T=618120 743000 1 0 $X=617830 $Y=738790
X584 6 5 ICV_47 $T=660120 633240 1 0 $X=659830 $Y=629030
X585 6 5 ICV_47 $T=660120 641080 0 0 $X=659830 $Y=640845
X586 6 5 ICV_47 $T=660120 688120 1 0 $X=659830 $Y=683910
X587 6 5 ICV_47 $T=660120 735160 1 0 $X=659830 $Y=730950
X588 6 5 ICV_47 $T=660120 743000 1 0 $X=659830 $Y=738790
X589 6 5 ICV_47 $T=702120 641080 1 0 $X=701830 $Y=636870
X590 6 5 ICV_47 $T=702120 680280 1 0 $X=701830 $Y=676070
X591 6 5 ICV_47 $T=702120 735160 1 0 $X=701830 $Y=730950
X592 5 6 DCAP32BWP7T $T=454040 648920 1 0 $X=453750 $Y=644710
X593 5 6 DCAP32BWP7T $T=461320 648920 0 0 $X=461030 $Y=648685
X594 5 6 DCAP32BWP7T $T=466920 688120 0 0 $X=466630 $Y=687885
X595 5 6 DCAP32BWP7T $T=469160 625400 1 0 $X=468870 $Y=621190
X596 5 6 DCAP32BWP7T $T=469160 719480 0 0 $X=468870 $Y=719245
X597 5 6 DCAP32BWP7T $T=473080 672440 1 0 $X=472790 $Y=668230
X598 5 6 DCAP32BWP7T $T=492120 633240 0 0 $X=491830 $Y=633005
X599 5 6 DCAP32BWP7T $T=492120 719480 1 0 $X=491830 $Y=715270
X600 5 6 DCAP32BWP7T $T=492120 743000 1 0 $X=491830 $Y=738790
X601 5 6 DCAP32BWP7T $T=515080 688120 0 0 $X=514790 $Y=687885
X602 5 6 DCAP32BWP7T $T=534120 601880 0 0 $X=533830 $Y=601645
X603 5 6 DCAP32BWP7T $T=534120 680280 0 0 $X=533830 $Y=680045
X604 5 6 DCAP32BWP7T $T=534120 727320 0 0 $X=533830 $Y=727085
X605 5 6 DCAP32BWP7T $T=534120 743000 1 0 $X=533830 $Y=738790
X606 5 6 DCAP32BWP7T $T=545320 695960 1 0 $X=545030 $Y=691750
X607 5 6 DCAP32BWP7T $T=548120 633240 0 0 $X=547830 $Y=633005
X608 5 6 DCAP32BWP7T $T=555960 609720 0 0 $X=555670 $Y=609485
X609 5 6 DCAP32BWP7T $T=555960 719480 1 0 $X=555670 $Y=715270
X610 5 6 DCAP32BWP7T $T=593480 672440 0 0 $X=593190 $Y=672205
X611 5 6 DCAP32BWP7T $T=598520 656760 0 0 $X=598230 $Y=656525
X612 5 6 DCAP32BWP7T $T=618120 601880 1 0 $X=617830 $Y=597670
X613 5 6 DCAP32BWP7T $T=618120 609720 1 0 $X=617830 $Y=605510
X614 5 6 DCAP32BWP7T $T=618120 641080 1 0 $X=617830 $Y=636870
X615 5 6 DCAP32BWP7T $T=618120 648920 0 0 $X=617830 $Y=648685
X616 5 6 DCAP32BWP7T $T=618120 656760 0 0 $X=617830 $Y=656525
X617 5 6 DCAP32BWP7T $T=618120 695960 1 0 $X=617830 $Y=691750
X618 5 6 DCAP32BWP7T $T=618120 719480 0 0 $X=617830 $Y=719245
X619 5 6 DCAP32BWP7T $T=660120 703800 1 0 $X=659830 $Y=699590
X620 5 6 DCAP32BWP7T $T=660120 711640 0 0 $X=659830 $Y=711405
X621 5 6 DCAP32BWP7T $T=660120 719480 1 0 $X=659830 $Y=715270
X622 5 6 DCAP32BWP7T $T=669640 672440 1 0 $X=669350 $Y=668230
X623 5 6 DCAP32BWP7T $T=682520 711640 1 0 $X=682230 $Y=707430
X624 5 6 DCAP32BWP7T $T=702120 656760 1 0 $X=701830 $Y=652550
X625 5 6 DCAP32BWP7T $T=709960 695960 1 0 $X=709670 $Y=691750
X626 5 6 DCAP32BWP7T $T=716120 672440 0 0 $X=715830 $Y=672205
X627 5 6 DCAP32BWP7T $T=719480 743000 1 0 $X=719190 $Y=738790
X628 5 6 DCAP32BWP7T $T=724520 633240 0 0 $X=724230 $Y=633005
X629 34 188 196 204 5 6 207 FA1D0BWP7T $T=456280 711640 1 0 $X=455990 $Y=707430
X630 7 192 202 205 5 6 206 FA1D0BWP7T $T=456280 719480 0 0 $X=455990 $Y=719245
X631 37 45 55 210 5 6 213 FA1D0BWP7T $T=459640 641080 0 0 $X=459350 $Y=640845
X632 38 48 183 58 5 6 214 FA1D0BWP7T $T=460200 656760 1 0 $X=459910 $Y=652550
X633 40 199 209 212 5 6 215 FA1D0BWP7T $T=460200 672440 1 0 $X=459910 $Y=668230
X634 208 61 216 227 5 6 230 FA1D0BWP7T $T=469720 727320 1 0 $X=469430 $Y=723110
X635 182 201 195 228 5 6 233 FA1D0BWP7T $T=470280 711640 1 0 $X=469990 $Y=707430
X636 205 66 204 209 5 6 240 FA1D0BWP7T $T=471960 695960 0 0 $X=471670 $Y=695725
X637 74 241 189 242 5 6 278 FA1D0BWP7T $T=492680 633240 1 0 $X=492390 $Y=629030
X638 280 228 207 255 5 6 248 FA1D0BWP7T $T=505560 680280 1 180 $X=492390 $Y=680045
X639 232 217 244 88 5 6 89 FA1D0BWP7T $T=493240 617560 1 0 $X=492950 $Y=613350
X640 279 275 261 260 5 6 257 FA1D0BWP7T $T=507240 735160 1 180 $X=494070 $Y=734925
X641 227 233 260 285 5 6 287 FA1D0BWP7T $T=497160 711640 1 0 $X=496870 $Y=707430
X642 219 269 206 280 5 6 289 FA1D0BWP7T $T=497160 719480 0 0 $X=496870 $Y=719245
X643 251 271 295 298 5 6 288 FA1D0BWP7T $T=503880 625400 0 0 $X=503590 $Y=625165
X644 259 284 248 299 5 6 319 FA1D0BWP7T $T=503880 664600 0 0 $X=503590 $Y=664365
X645 184 264 263 306 5 6 309 FA1D0BWP7T $T=506680 641080 1 0 $X=506390 $Y=636870
X646 312 304 252 269 5 6 286 FA1D0BWP7T $T=521800 735160 0 180 $X=508630 $Y=730950
X647 286 62 311 315 5 6 317 FA1D0BWP7T $T=510600 703800 0 0 $X=510310 $Y=703565
X648 253 303 282 320 5 6 281 FA1D0BWP7T $T=512840 601880 0 0 $X=512550 $Y=601645
X649 267 254 220 321 5 6 326 FA1D0BWP7T $T=512840 656760 1 0 $X=512550 $Y=652550
X650 298 310 320 327 5 6 334 FA1D0BWP7T $T=515640 633240 1 0 $X=515350 $Y=629030
X651 245 306 322 308 5 6 335 FA1D0BWP7T $T=515640 641080 0 0 $X=515350 $Y=640845
X652 315 285 289 284 5 6 301 FA1D0BWP7T $T=528520 680280 1 180 $X=515350 $Y=680045
X653 326 346 357 361 5 6 358 FA1D0BWP7T $T=535800 641080 0 0 $X=535510 $Y=640845
X654 283 101 268 364 5 6 366 FA1D0BWP7T $T=539160 656760 0 0 $X=538870 $Y=656525
X655 362 321 366 382 5 6 383 FA1D0BWP7T $T=547560 672440 1 0 $X=547270 $Y=668230
X656 386 378 355 363 5 6 310 FA1D0BWP7T $T=560440 688120 0 180 $X=547270 $Y=683910
X657 361 327 383 387 5 6 296 FA1D0BWP7T $T=549240 641080 0 0 $X=548950 $Y=640845
X658 335 379 400 403 5 6 407 FA1D0BWP7T $T=557640 648920 0 0 $X=557350 $Y=648685
X659 364 309 397 400 5 6 409 FA1D0BWP7T $T=557640 664600 0 0 $X=557350 $Y=664365
X660 377 388 365 397 5 6 408 FA1D0BWP7T $T=557640 680280 0 0 $X=557350 $Y=680045
X661 411 387 418 420 5 6 373 FA1D0BWP7T $T=576680 609720 0 0 $X=576390 $Y=609485
X662 382 363 408 415 5 6 418 FA1D0BWP7T $T=576680 656760 0 0 $X=576390 $Y=656525
X663 121 116 113 414 5 6 112 FA1D0BWP7T $T=593480 601880 0 180 $X=580310 $Y=597670
X664 118 414 126 422 5 6 437 FA1D0BWP7T $T=592920 609720 1 0 $X=592630 $Y=605510
X665 453 137 437 459 5 6 133 FA1D0BWP7T $T=632680 601880 1 180 $X=619510 $Y=601645
X666 19 6 5 180 INVD1BWP7T $T=452360 711640 1 180 $X=450390 $Y=711405
X667 15 6 5 20 INVD1BWP7T $T=450680 727320 1 0 $X=450390 $Y=723110
X668 8 6 5 24 INVD1BWP7T $T=463560 695960 1 180 $X=461590 $Y=695725
X669 246 6 5 32 INVD1BWP7T $T=486520 735160 1 180 $X=484550 $Y=734925
X670 272 6 5 266 INVD1BWP7T $T=502200 641080 1 180 $X=500230 $Y=640845
X671 292 6 5 92 INVD1BWP7T $T=511720 743000 0 180 $X=509750 $Y=738790
X672 300 6 5 46 INVD1BWP7T $T=516760 719480 1 180 $X=514790 $Y=719245
X673 374 6 5 53 INVD1BWP7T $T=558760 735160 1 180 $X=556790 $Y=734925
X674 371 6 5 28 INVD1BWP7T $T=562680 695960 1 180 $X=560710 $Y=695725
X675 384 6 5 256 INVD1BWP7T $T=581160 688120 0 180 $X=579190 $Y=683910
X676 404 6 5 273 INVD1BWP7T $T=582840 695960 1 180 $X=580870 $Y=695725
X677 128 6 5 229 INVD1BWP7T $T=607480 672440 0 180 $X=605510 $Y=668230
X678 142 6 5 134 INVD1BWP7T $T=638840 609720 0 180 $X=636870 $Y=605510
X679 141 6 5 80 INVD1BWP7T $T=639960 601880 0 180 $X=637990 $Y=597670
X827 237 6 218 18 5 ND2D1BWP7T $T=484840 735160 1 180 $X=482310 $Y=734925
X828 246 6 236 18 5 ND2D1BWP7T $T=486520 735160 0 180 $X=483990 $Y=730950
X829 258 6 250 8 5 ND2D1BWP7T $T=494920 719480 1 180 $X=492390 $Y=719245
X830 83 6 84 85 5 ND2D1BWP7T $T=494920 601880 0 0 $X=494630 $Y=601645
X831 29 6 291 93 5 ND2D1BWP7T $T=509480 695960 0 0 $X=509190 $Y=695725
X832 297 6 307 18 5 ND2D1BWP7T $T=516760 719480 0 0 $X=516470 $Y=719245
X833 337 6 329 292 5 ND2D1BWP7T $T=528520 743000 0 180 $X=525990 $Y=738790
X834 99 6 341 85 5 ND2D1BWP7T $T=539720 633240 0 0 $X=539430 $Y=633005
X835 100 6 348 98 5 ND2D1BWP7T $T=540280 601880 1 0 $X=539990 $Y=597670
X836 237 6 354 300 5 ND2D1BWP7T $T=545320 727320 0 180 $X=542790 $Y=723110
X837 77 6 360 272 5 ND2D1BWP7T $T=545880 633240 0 0 $X=545590 $Y=633005
X838 246 6 356 374 5 ND2D1BWP7T $T=557080 735160 1 180 $X=554550 $Y=734925
X839 15 6 345 347 5 ND2D1BWP7T $T=570520 703800 0 180 $X=567990 $Y=699590
X840 384 6 376 107 5 ND2D1BWP7T $T=577800 641080 1 0 $X=577510 $Y=636870
X841 19 6 352 72 5 ND2D1BWP7T $T=580040 672440 0 0 $X=579750 $Y=672205
X842 371 6 396 123 5 ND2D1BWP7T $T=593480 617560 0 0 $X=593190 $Y=617325
X843 404 6 385 128 5 ND2D1BWP7T $T=629880 633240 0 180 $X=627350 $Y=629030
X844 130 6 140 141 5 ND2D1BWP7T $T=636040 601880 1 0 $X=635750 $Y=597670
X845 151 6 457 149 5 ND2D1BWP7T $T=653400 609720 1 180 $X=650870 $Y=609485
X846 168 6 143 163 5 ND2D1BWP7T $T=690360 609720 0 180 $X=687830 $Y=605510
X847 151 6 440 163 5 ND2D1BWP7T $T=688120 656760 1 0 $X=687830 $Y=652550
X848 151 6 456 167 5 ND2D1BWP7T $T=688680 648920 1 0 $X=688390 $Y=644710
X849 553 6 405 166 5 ND2D1BWP7T $T=690920 672440 1 180 $X=688390 $Y=672205
X850 151 6 431 170 5 ND2D1BWP7T $T=690920 648920 1 0 $X=690630 $Y=644710
X880 16 6 5 186 INVD0BWP7T $T=450680 703800 0 0 $X=450390 $Y=703565
X881 31 6 5 33 INVD0BWP7T $T=454040 735160 1 0 $X=453750 $Y=730950
X882 200 6 5 199 INVD0BWP7T $T=465240 695960 1 180 $X=463270 $Y=695725
X883 242 6 5 244 INVD0BWP7T $T=484840 617560 1 0 $X=484550 $Y=613350
X884 238 6 5 245 INVD0BWP7T $T=484840 617560 0 0 $X=484550 $Y=617325
X885 213 6 5 222 INVD0BWP7T $T=486520 641080 0 180 $X=484550 $Y=636870
X886 313 6 5 379 INVD0BWP7T $T=555400 656760 1 0 $X=555110 $Y=652550
X887 11 197 185 49 6 5 OAI21D0BWP7T $T=468600 625400 1 180 $X=465510 $Y=625165
X888 203 232 73 238 6 5 OAI21D0BWP7T $T=482040 617560 0 0 $X=481750 $Y=617325
X889 240 249 255 215 6 5 OAI21D0BWP7T $T=492680 703800 0 0 $X=492390 $Y=703565
X890 96 402 405 393 6 5 OAI21D0BWP7T $T=567720 727320 1 0 $X=567430 $Y=723110
X891 96 412 413 342 6 5 OAI21D0BWP7T $T=577800 735160 0 0 $X=577510 $Y=734925
X892 413 445 106 417 6 5 OAI21D0BWP7T $T=581720 727320 0 0 $X=581430 $Y=727085
X893 409 427 415 407 6 5 OAI21D0BWP7T $T=582280 672440 1 0 $X=581990 $Y=668230
X894 117 424 422 115 6 5 OAI21D0BWP7T $T=590680 633240 0 180 $X=587590 $Y=629030
X895 96 429 431 421 6 5 OAI21D0BWP7T $T=599640 695960 1 180 $X=596550 $Y=695725
X896 405 435 106 450 6 5 OAI21D0BWP7T $T=601880 719480 1 0 $X=601590 $Y=715270
X897 96 436 440 443 6 5 OAI21D0BWP7T $T=605800 680280 1 0 $X=605510 $Y=676070
X898 324 441 106 438 6 5 OAI21D0BWP7T $T=608600 727320 0 180 $X=605510 $Y=723110
X899 431 451 106 454 6 5 OAI21D0BWP7T $T=609720 695960 0 0 $X=609430 $Y=695725
X900 96 448 457 460 6 5 OAI21D0BWP7T $T=618680 648920 1 0 $X=618390 $Y=644710
X901 96 432 456 425 6 5 OAI21D0BWP7T $T=621480 688120 0 180 $X=618390 $Y=683910
X902 135 461 413 464 6 5 OAI21D0BWP7T $T=620360 711640 0 0 $X=620070 $Y=711405
X903 457 458 106 465 6 5 OAI21D0BWP7T $T=627080 656760 0 180 $X=623990 $Y=652550
X904 135 484 323 466 6 5 OAI21D0BWP7T $T=624840 727320 0 0 $X=624550 $Y=727085
X905 440 470 106 472 6 5 OAI21D0BWP7T $T=634360 680280 1 180 $X=631270 $Y=680045
X906 456 468 106 480 6 5 OAI21D0BWP7T $T=633800 672440 1 0 $X=633510 $Y=668230
X907 135 485 324 477 6 5 OAI21D0BWP7T $T=641080 727320 0 180 $X=637990 $Y=723110
X908 135 486 457 483 6 5 OAI21D0BWP7T $T=641640 648920 1 180 $X=638550 $Y=648685
X909 135 488 431 500 6 5 OAI21D0BWP7T $T=641080 703800 1 0 $X=640790 $Y=699590
X910 135 491 405 473 6 5 OAI21D0BWP7T $T=643880 719480 0 180 $X=640790 $Y=715270
X911 457 493 146 489 6 5 OAI21D0BWP7T $T=645560 641080 0 180 $X=642470 $Y=636870
X912 143 496 147 492 6 5 OAI21D0BWP7T $T=646680 617560 1 180 $X=643590 $Y=617325
X913 135 474 456 498 6 5 OAI21D0BWP7T $T=644440 664600 1 0 $X=644150 $Y=660390
X914 324 494 146 499 6 5 OAI21D0BWP7T $T=644440 719480 0 0 $X=644150 $Y=719245
X915 456 505 146 536 6 5 OAI21D0BWP7T $T=650600 656760 0 0 $X=650310 $Y=656525
X916 135 504 440 501 6 5 OAI21D0BWP7T $T=653960 680280 1 180 $X=650870 $Y=680045
X917 413 508 146 515 6 5 OAI21D0BWP7T $T=651160 719480 0 0 $X=650870 $Y=719245
X918 150 511 457 513 6 5 OAI21D0BWP7T $T=651720 633240 0 0 $X=651430 $Y=633005
X919 405 510 146 514 6 5 OAI21D0BWP7T $T=651720 703800 0 0 $X=651430 $Y=703565
X920 152 495 143 516 6 5 OAI21D0BWP7T $T=660680 609720 1 0 $X=660390 $Y=605510
X921 431 529 146 518 6 5 OAI21D0BWP7T $T=660680 695960 0 0 $X=660390 $Y=695725
X922 154 523 457 525 6 5 OAI21D0BWP7T $T=664040 641080 1 0 $X=663750 $Y=636870
X923 156 517 143 526 6 5 OAI21D0BWP7T $T=671880 625400 0 180 $X=668790 $Y=621190
X924 440 519 146 537 6 5 OAI21D0BWP7T $T=672440 680280 1 0 $X=672150 $Y=676070
X925 158 538 143 532 6 5 OAI21D0BWP7T $T=676920 609720 1 180 $X=673830 $Y=609485
X926 143 533 155 522 6 5 OAI21D0BWP7T $T=679160 601880 1 180 $X=676070 $Y=601645
X927 150 542 324 531 6 5 OAI21D0BWP7T $T=679720 719480 0 0 $X=679430 $Y=719245
X928 324 534 154 546 6 5 OAI21D0BWP7T $T=681960 719480 1 0 $X=681670 $Y=715270
X929 152 543 162 552 6 5 OAI21D0BWP7T $T=684760 609720 0 0 $X=684470 $Y=609485
X930 150 549 405 556 6 5 OAI21D0BWP7T $T=687000 703800 1 0 $X=686710 $Y=699590
X931 456 545 154 561 6 5 OAI21D0BWP7T $T=687560 648920 0 0 $X=687270 $Y=648685
X932 150 548 456 560 6 5 OAI21D0BWP7T $T=688120 688120 0 0 $X=687830 $Y=687885
X933 169 551 155 559 6 5 OAI21D0BWP7T $T=693160 601880 1 180 $X=690070 $Y=601645
X934 150 566 413 564 6 5 OAI21D0BWP7T $T=694840 719480 1 180 $X=691750 $Y=719245
X935 152 563 169 565 6 5 OAI21D0BWP7T $T=696520 633240 1 180 $X=693430 $Y=633005
X936 323 557 146 554 6 5 OAI21D0BWP7T $T=702680 735160 0 0 $X=702390 $Y=734925
X937 440 580 154 575 6 5 OAI21D0BWP7T $T=708840 664600 0 180 $X=705750 $Y=660390
X938 323 579 154 598 6 5 OAI21D0BWP7T $T=706600 711640 0 0 $X=706310 $Y=711405
X939 150 581 431 585 6 5 OAI21D0BWP7T $T=707160 695960 1 0 $X=706870 $Y=691750
X940 158 584 169 574 6 5 OAI21D0BWP7T $T=710520 625400 1 180 $X=707430 $Y=625165
X941 158 583 162 588 6 5 OAI21D0BWP7T $T=708280 617560 1 0 $X=707990 $Y=613350
X942 405 586 154 589 6 5 OAI21D0BWP7T $T=708840 695960 0 0 $X=708550 $Y=695725
X943 150 590 440 568 6 5 OAI21D0BWP7T $T=712760 664600 1 180 $X=709670 $Y=664365
X944 156 595 169 594 6 5 OAI21D0BWP7T $T=718360 625400 1 180 $X=715270 $Y=625165
X945 150 582 323 578 6 5 OAI21D0BWP7T $T=716680 743000 1 0 $X=716390 $Y=738790
X946 156 604 162 601 6 5 OAI21D0BWP7T $T=725640 625400 1 180 $X=722550 $Y=625165
X947 169 602 147 600 6 5 OAI21D0BWP7T $T=727320 617560 0 180 $X=724230 $Y=613350
X948 413 606 154 610 6 5 OAI21D0BWP7T $T=733480 735160 1 180 $X=730390 $Y=734925
X949 162 621 147 614 6 5 OAI21D0BWP7T $T=735720 625400 1 0 $X=735430 $Y=621190
X950 431 620 154 605 6 5 OAI21D0BWP7T $T=738520 688120 1 180 $X=735430 $Y=687885
X1001 274 6 272 85 5 276 ND3D0BWP7T $T=502200 641080 0 0 $X=501910 $Y=640845
X1002 73 6 83 77 5 238 ND3D0BWP7T $T=512840 633240 0 0 $X=512550 $Y=633005
X1003 60 6 347 18 5 359 ND3D0BWP7T $T=557640 727320 1 0 $X=557350 $Y=723110
X1004 6 5 DCAP16BWP7T $T=450120 641080 0 0 $X=449830 $Y=640845
X1005 6 5 DCAP16BWP7T $T=450120 656760 1 0 $X=449830 $Y=652550
X1006 6 5 DCAP16BWP7T $T=456840 727320 1 0 $X=456550 $Y=723110
X1007 6 5 DCAP16BWP7T $T=461320 664600 1 0 $X=461030 $Y=660390
X1008 6 5 DCAP16BWP7T $T=468040 601880 0 0 $X=467750 $Y=601645
X1009 6 5 DCAP16BWP7T $T=479240 688120 1 0 $X=478950 $Y=683910
X1010 6 5 DCAP16BWP7T $T=480360 601880 0 0 $X=480070 $Y=601645
X1011 6 5 DCAP16BWP7T $T=492120 601880 1 0 $X=491830 $Y=597670
X1012 6 5 DCAP16BWP7T $T=492120 625400 0 0 $X=491830 $Y=625165
X1013 6 5 DCAP16BWP7T $T=492120 680280 1 0 $X=491830 $Y=676070
X1014 6 5 DCAP16BWP7T $T=492120 688120 0 0 $X=491830 $Y=687885
X1015 6 5 DCAP16BWP7T $T=494920 695960 0 0 $X=494630 $Y=695725
X1016 6 5 DCAP16BWP7T $T=495480 703800 0 0 $X=495190 $Y=703565
X1017 6 5 DCAP16BWP7T $T=502760 672440 1 0 $X=502470 $Y=668230
X1018 6 5 DCAP16BWP7T $T=503880 695960 1 0 $X=503590 $Y=691750
X1019 6 5 DCAP16BWP7T $T=505560 680280 0 0 $X=505270 $Y=680045
X1020 6 5 DCAP16BWP7T $T=511720 743000 1 0 $X=511430 $Y=738790
X1021 6 5 DCAP16BWP7T $T=515080 727320 1 0 $X=514790 $Y=723110
X1022 6 5 DCAP16BWP7T $T=523480 703800 0 0 $X=523190 $Y=703565
X1023 6 5 DCAP16BWP7T $T=534120 617560 1 0 $X=533830 $Y=613350
X1024 6 5 DCAP16BWP7T $T=534120 695960 1 0 $X=533830 $Y=691750
X1025 6 5 DCAP16BWP7T $T=534120 727320 1 0 $X=533830 $Y=723110
X1026 6 5 DCAP16BWP7T $T=555400 743000 1 0 $X=555110 $Y=738790
X1027 6 5 DCAP16BWP7T $T=555960 727320 0 0 $X=555670 $Y=727085
X1028 6 5 DCAP16BWP7T $T=562120 641080 0 0 $X=561830 $Y=640845
X1029 6 5 DCAP16BWP7T $T=564360 719480 0 0 $X=564070 $Y=719245
X1030 6 5 DCAP16BWP7T $T=576120 703800 1 0 $X=575830 $Y=699590
X1031 6 5 DCAP16BWP7T $T=576120 711640 0 0 $X=575830 $Y=711405
X1032 6 5 DCAP16BWP7T $T=578920 633240 1 0 $X=578630 $Y=629030
X1033 6 5 DCAP16BWP7T $T=599640 695960 0 0 $X=599350 $Y=695725
X1034 6 5 DCAP16BWP7T $T=604680 719480 1 0 $X=604390 $Y=715270
X1035 6 5 DCAP16BWP7T $T=606360 641080 0 0 $X=606070 $Y=640845
X1036 6 5 DCAP16BWP7T $T=607480 672440 1 0 $X=607190 $Y=668230
X1037 6 5 DCAP16BWP7T $T=607480 680280 0 0 $X=607190 $Y=680045
X1038 6 5 DCAP16BWP7T $T=618120 695960 0 0 $X=617830 $Y=695725
X1039 6 5 DCAP16BWP7T $T=629320 703800 1 0 $X=629030 $Y=699590
X1040 6 5 DCAP16BWP7T $T=632120 680280 1 0 $X=631830 $Y=676070
X1041 6 5 DCAP16BWP7T $T=638840 633240 0 0 $X=638550 $Y=633005
X1042 6 5 DCAP16BWP7T $T=647240 664600 1 0 $X=646950 $Y=660390
X1043 6 5 DCAP16BWP7T $T=647800 617560 1 0 $X=647510 $Y=613350
X1044 6 5 DCAP16BWP7T $T=647800 633240 1 0 $X=647510 $Y=629030
X1045 6 5 DCAP16BWP7T $T=649480 680280 1 0 $X=649190 $Y=676070
X1046 6 5 DCAP16BWP7T $T=660120 609720 0 0 $X=659830 $Y=609485
X1047 6 5 DCAP16BWP7T $T=660120 625400 1 0 $X=659830 $Y=621190
X1048 6 5 DCAP16BWP7T $T=660120 680280 1 0 $X=659830 $Y=676070
X1049 6 5 DCAP16BWP7T $T=669080 617560 1 0 $X=668790 $Y=613350
X1050 6 5 DCAP16BWP7T $T=679160 601880 0 0 $X=678870 $Y=601645
X1051 6 5 DCAP16BWP7T $T=682520 719480 0 0 $X=682230 $Y=719245
X1052 6 5 DCAP16BWP7T $T=688680 719480 1 0 $X=688390 $Y=715270
X1053 6 5 DCAP16BWP7T $T=689240 601880 1 0 $X=688950 $Y=597670
X1054 6 5 DCAP16BWP7T $T=689800 703800 1 0 $X=689510 $Y=699590
X1055 6 5 DCAP16BWP7T $T=690360 609720 1 0 $X=690070 $Y=605510
X1056 6 5 DCAP16BWP7T $T=690360 648920 0 0 $X=690070 $Y=648685
X1057 6 5 DCAP16BWP7T $T=690920 672440 0 0 $X=690630 $Y=672205
X1058 6 5 DCAP16BWP7T $T=690920 688120 0 0 $X=690630 $Y=687885
X1059 6 5 DCAP16BWP7T $T=692040 664600 0 0 $X=691750 $Y=664365
X1060 6 5 DCAP16BWP7T $T=702120 672440 1 0 $X=701830 $Y=668230
X1061 6 5 DCAP16BWP7T $T=702120 680280 0 0 $X=701830 $Y=680045
X1062 6 5 DCAP16BWP7T $T=702120 688120 0 0 $X=701830 $Y=687885
X1063 6 5 DCAP16BWP7T $T=716120 727320 1 0 $X=715830 $Y=723110
X1064 6 5 DCAP16BWP7T $T=723400 719480 1 0 $X=723110 $Y=715270
X1110 21 6 180 9 34 5 NR3D1BWP7T $T=450680 719480 1 0 $X=450390 $Y=715270
X1111 21 6 32 186 182 5 NR3D1BWP7T $T=452360 727320 1 0 $X=452070 $Y=723110
X1112 224 6 187 76 74 5 NR3D1BWP7T $T=484280 625400 1 180 $X=479510 $Y=625165
X1113 222 64 6 5 214 200 MAOI222D1BWP7T $T=478680 641080 1 180 $X=473910 $Y=640845
X1114 95 308 6 5 278 313 MAOI222D1BWP7T $T=516760 617560 0 0 $X=516470 $Y=617325
X1115 33 218 6 62 219 5 AOI21D1BWP7T $T=478120 735160 1 180 $X=474470 $Y=734925
X1116 29 14 5 6 INVD2BWP7T $T=453480 695960 1 180 $X=450950 $Y=695725
X1117 18 21 5 6 INVD2BWP7T $T=451240 735160 0 0 $X=450950 $Y=734925
X1118 77 23 5 6 INVD2BWP7T $T=484840 633240 0 180 $X=482310 $Y=629030
X1119 83 187 5 6 INVD2BWP7T $T=502760 601880 0 0 $X=502470 $Y=601645
X1120 103 179 5 6 INVD2BWP7T $T=545880 617560 1 0 $X=545590 $Y=613350
X1121 337 44 5 6 INVD2BWP7T $T=555400 743000 0 180 $X=552870 $Y=738790
X1122 85 224 5 6 INVD2BWP7T $T=580600 695960 0 180 $X=578070 $Y=691750
X1195 36 43 6 5 27 DFQD0BWP7T $T=464120 601880 0 180 $X=453190 $Y=597670
X1196 36 42 6 5 54 DFQD0BWP7T $T=458520 625400 1 0 $X=458230 $Y=621190
X1197 36 52 6 5 50 DFQD0BWP7T $T=465800 609720 1 0 $X=465510 $Y=605510
X1198 36 94 6 5 258 DFQD0BWP7T $T=515080 688120 1 180 $X=504150 $Y=687885
X1199 36 97 6 5 297 DFQD0BWP7T $T=526840 695960 0 180 $X=515910 $Y=691750
X1200 36 349 6 5 305 DFQD0BWP7T $T=545320 609720 1 180 $X=534390 $Y=609485
X1201 102 330 6 5 347 DFQD0BWP7T $T=550360 695960 1 180 $X=539430 $Y=695725
X1202 36 368 6 5 272 DFQD0BWP7T $T=555960 609720 1 180 $X=545030 $Y=609485
X1203 102 367 6 5 337 DFQD0BWP7T $T=555960 711640 0 180 $X=545030 $Y=707430
X1204 102 353 6 5 380 DFQD0BWP7T $T=567720 711640 0 180 $X=556790 $Y=707430
X1205 36 391 6 5 375 DFQD0BWP7T $T=568280 617560 0 180 $X=557350 $Y=613350
X1206 102 395 6 5 384 DFQD0BWP7T $T=569960 633240 0 180 $X=559030 $Y=629030
X1207 102 406 6 5 410 DFQD0BWP7T $T=587320 625400 1 180 $X=576390 $Y=625165
X1208 102 416 6 5 262 DFQD0BWP7T $T=587320 641080 1 180 $X=576390 $Y=640845
X1209 102 122 6 5 114 DFQD0BWP7T $T=597960 625400 1 180 $X=587030 $Y=625165
X1210 102 430 6 5 302 DFQD0BWP7T $T=600760 664600 1 180 $X=589830 $Y=664365
X1211 102 394 6 5 325 DFQD0BWP7T $T=593480 735160 0 0 $X=593190 $Y=734925
X1212 102 439 6 5 434 DFQD0BWP7T $T=610280 625400 1 180 $X=599350 $Y=625165
X1213 102 446 6 5 125 DFQD0BWP7T $T=612520 641080 0 180 $X=601590 $Y=636870
X1214 102 447 6 5 274 DFQD0BWP7T $T=612520 656760 0 180 $X=601590 $Y=652550
X1215 102 435 6 5 399 DFQD0BWP7T $T=601880 703800 0 0 $X=601590 $Y=703565
X1216 102 445 6 5 340 DFQD0BWP7T $T=612520 735160 0 180 $X=601590 $Y=730950
X1217 102 458 6 5 462 DFQD0BWP7T $T=618680 664600 0 0 $X=618390 $Y=664365
X1218 102 451 6 5 419 DFQD0BWP7T $T=629320 703800 0 180 $X=618390 $Y=699590
X1219 102 441 6 5 398 DFQD0BWP7T $T=631000 735160 1 180 $X=620070 $Y=734925
X1220 102 468 6 5 426 DFQD0BWP7T $T=632120 680280 0 180 $X=621190 $Y=676070
X1221 102 470 6 5 444 DFQD0BWP7T $T=633240 688120 1 180 $X=622310 $Y=687885
X1222 102 461 6 5 442 DFQD0BWP7T $T=639400 711640 0 180 $X=628470 $Y=707430
X1223 102 474 6 5 487 DFQD0BWP7T $T=631000 664600 0 0 $X=630710 $Y=664365
X1224 102 476 6 5 478 DFQD0BWP7T $T=632120 625400 0 0 $X=631830 $Y=625165
X1225 102 484 6 5 401 DFQD0BWP7T $T=643320 735160 1 180 $X=632390 $Y=734925
X1226 102 486 6 5 471 DFQD0BWP7T $T=643880 656760 0 180 $X=632950 $Y=652550
X1227 102 488 6 5 479 DFQD0BWP7T $T=646680 695960 0 180 $X=635750 $Y=691750
X1228 102 491 6 5 455 DFQD0BWP7T $T=651720 711640 0 180 $X=640790 $Y=707430
X1229 102 495 6 5 512 DFQD0BWP7T $T=643320 601880 0 0 $X=643030 $Y=601645
X1230 102 504 6 5 490 DFQD0BWP7T $T=653960 672440 0 180 $X=643030 $Y=668230
X1231 102 496 6 5 497 DFQD0BWP7T $T=643880 625400 0 0 $X=643590 $Y=625165
X1232 102 493 6 5 482 DFQD0BWP7T $T=654520 641080 1 180 $X=643590 $Y=640845
X1233 102 485 6 5 463 DFQD0BWP7T $T=654520 735160 1 180 $X=643590 $Y=734925
X1234 102 517 6 5 524 DFQD0BWP7T $T=660680 625400 0 0 $X=660390 $Y=625165
X1235 102 505 6 5 503 DFQD0BWP7T $T=671320 664600 1 180 $X=660390 $Y=664365
X1236 102 510 6 5 475 DFQD0BWP7T $T=671320 711640 0 180 $X=660390 $Y=707430
X1237 102 494 6 5 481 DFQD0BWP7T $T=660680 735160 0 0 $X=660390 $Y=734925
X1238 102 519 6 5 506 DFQD0BWP7T $T=661800 680280 0 0 $X=661510 $Y=680045
X1239 102 529 6 5 502 DFQD0BWP7T $T=672440 695960 0 180 $X=661510 $Y=691750
X1240 102 511 6 5 509 DFQD0BWP7T $T=673000 656760 0 180 $X=662070 $Y=652550
X1241 102 533 6 5 153 DFQD0BWP7T $T=676360 601880 0 180 $X=665430 $Y=597670
X1242 102 508 6 5 467 DFQD0BWP7T $T=679160 727320 0 180 $X=668230 $Y=723110
X1243 102 542 6 5 507 DFQD0BWP7T $T=681960 735160 1 180 $X=671030 $Y=734925
X1244 102 534 6 5 527 DFQD0BWP7T $T=671880 711640 1 0 $X=671590 $Y=707430
X1245 102 538 6 5 520 DFQD0BWP7T $T=683080 625400 1 180 $X=672150 $Y=625165
X1246 102 523 6 5 528 DFQD0BWP7T $T=685880 656760 0 180 $X=674950 $Y=652550
X1247 102 535 6 5 530 DFQD0BWP7T $T=677480 641080 1 0 $X=677190 $Y=636870
X1248 102 551 6 5 161 DFQD0BWP7T $T=689240 601880 0 180 $X=678310 $Y=597670
X1249 102 543 6 5 165 DFQD0BWP7T $T=678600 617560 1 0 $X=678310 $Y=613350
X1250 102 548 6 5 540 DFQD0BWP7T $T=689240 680280 1 180 $X=678310 $Y=680045
X1251 102 549 6 5 541 DFQD0BWP7T $T=689240 695960 0 180 $X=678310 $Y=691750
X1252 102 545 6 5 562 DFQD0BWP7T $T=681400 664600 0 0 $X=681110 $Y=664365
X1253 102 557 6 5 469 DFQD0BWP7T $T=693160 735160 1 180 $X=682230 $Y=734925
X1254 102 550 6 5 555 DFQD0BWP7T $T=683640 703800 0 0 $X=683350 $Y=703565
X1255 102 563 6 5 547 DFQD0BWP7T $T=695400 625400 1 180 $X=684470 $Y=625165
X1256 102 584 6 5 572 DFQD0BWP7T $T=713320 633240 1 180 $X=702390 $Y=633005
X1257 102 583 6 5 573 DFQD0BWP7T $T=714440 609720 0 180 $X=703510 $Y=605510
X1258 102 581 6 5 539 DFQD0BWP7T $T=715000 688120 0 180 $X=704070 $Y=683910
X1259 102 576 6 5 567 DFQD0BWP7T $T=715560 648920 0 180 $X=704630 $Y=644710
X1260 102 590 6 5 544 DFQD0BWP7T $T=716120 672440 1 180 $X=705190 $Y=672205
X1261 102 566 6 5 521 DFQD0BWP7T $T=716120 727320 0 180 $X=705190 $Y=723110
X1262 102 582 6 5 558 DFQD0BWP7T $T=706600 735160 0 0 $X=706310 $Y=734925
X1263 102 579 6 5 587 DFQD0BWP7T $T=707160 711640 1 0 $X=706870 $Y=707430
X1264 102 595 6 5 591 DFQD0BWP7T $T=724520 633240 1 180 $X=713590 $Y=633005
X1265 102 586 6 5 569 DFQD0BWP7T $T=724520 695960 1 180 $X=713590 $Y=695725
X1266 102 602 6 5 596 DFQD0BWP7T $T=727320 609720 0 180 $X=716390 $Y=605510
X1267 102 604 6 5 592 DFQD0BWP7T $T=727880 648920 0 180 $X=716950 $Y=644710
X1268 102 580 6 5 571 DFQD0BWP7T $T=727880 672440 0 180 $X=716950 $Y=668230
X1269 102 606 6 5 570 DFQD0BWP7T $T=729000 727320 1 180 $X=718070 $Y=727085
X1270 102 593 6 5 577 DFQD0BWP7T $T=729560 656760 1 180 $X=718630 $Y=656525
X1271 102 617 6 5 603 DFQD0BWP7T $T=738520 601880 1 180 $X=727590 $Y=601645
X1272 102 621 6 5 607 DFQD0BWP7T $T=738520 633240 0 180 $X=727590 $Y=629030
X1273 102 618 6 5 612 DFQD0BWP7T $T=738520 641080 1 180 $X=727590 $Y=640845
X1274 102 619 6 5 608 DFQD0BWP7T $T=738520 672440 0 180 $X=727590 $Y=668230
X1275 102 620 6 5 597 DFQD0BWP7T $T=738520 680280 1 180 $X=727590 $Y=680045
X1276 102 609 6 5 599 DFQD0BWP7T $T=738520 695960 1 180 $X=727590 $Y=695725
X1277 102 615 6 5 611 DFQD0BWP7T $T=738520 711640 0 180 $X=727590 $Y=707430
X1278 102 616 6 5 613 DFQD0BWP7T $T=738520 727320 0 180 $X=727590 $Y=723110
X1279 236 188 186 182 6 5 AOI21D0BWP7T $T=453480 703800 0 180 $X=450390 $Y=699590
X1280 297 8 6 5 275 AN2D1BWP7T $T=515080 719480 1 180 $X=511990 $Y=719245
X1281 99 98 6 5 303 AN2D1BWP7T $T=537480 601880 0 180 $X=534390 $Y=597670
X1282 347 8 6 5 312 AN2D1BWP7T $T=542520 719480 1 180 $X=539430 $Y=719245
X1283 347 18 6 5 369 AN2D1BWP7T $T=556520 727320 0 180 $X=553430 $Y=723110
X1284 308 278 89 5 6 333 XOR3D0BWP7T $T=519000 617560 1 0 $X=518710 $Y=613350
X1285 17 30 35 5 6 41 XNR3D0BWP7T $T=450680 625400 0 0 $X=450390 $Y=625165
X1286 56 67 211 5 6 59 XNR3D0BWP7T $T=481480 617560 0 180 $X=471670 $Y=613350
X1287 240 215 255 5 6 270 XNR3D0BWP7T $T=492680 664600 0 0 $X=492390 $Y=664365
X1288 409 407 415 5 6 428 XNR3D0BWP7T $T=587320 641080 0 0 $X=587030 $Y=640845
X1289 117 115 422 5 6 452 XNR3D0BWP7T $T=601880 617560 0 0 $X=601590 $Y=617325
X1290 240 255 6 259 249 5 IOA21D0BWP7T $T=492680 711640 1 0 $X=492390 $Y=707430
X1291 409 415 6 411 427 5 IOA21D0BWP7T $T=598520 656760 1 180 $X=594870 $Y=656525
X1292 117 422 6 453 424 5 IOA21D0BWP7T $T=609160 609720 1 0 $X=608870 $Y=605510
X1293 290 91 212 51 6 5 194 AO22D0BWP7T $T=510600 656760 0 180 $X=505830 $Y=652550
X1294 274 91 299 51 6 5 225 AO22D0BWP7T $T=539160 656760 1 180 $X=534390 $Y=656525
X1295 125 91 420 51 6 5 447 AO22D0BWP7T $T=618680 633240 1 0 $X=618390 $Y=629030
X1296 114 91 403 51 6 5 433 AO22D0BWP7T $T=623160 633240 1 0 $X=622870 $Y=629030
X1297 145 91 459 51 6 5 446 AO22D0BWP7T $T=642200 609720 1 180 $X=637430 $Y=609485
X1298 56 211 57 217 6 5 MAOI222D2BWP7T $T=469160 625400 0 0 $X=468870 $Y=625165
X1299 36 190 6 5 11 DFQD1BWP7T $T=461320 633240 1 180 $X=450390 $Y=633005
X1300 36 193 6 5 12 DFQD1BWP7T $T=461320 648920 1 180 $X=450390 $Y=648685
X1301 36 191 6 5 13 DFQD1BWP7T $T=461320 664600 0 180 $X=450390 $Y=660390
X1302 36 39 6 5 25 DFQD1BWP7T $T=463560 609720 1 180 $X=452630 $Y=609485
X1303 36 194 6 5 16 DFQD1BWP7T $T=463560 680280 0 180 $X=452630 $Y=676070
X1304 36 198 6 5 31 DFQD1BWP7T $T=466920 688120 1 180 $X=455990 $Y=687885
X1305 36 181 6 5 29 DFQD1BWP7T $T=479240 688120 0 180 $X=468310 $Y=683910
X1306 36 234 6 5 65 DFQD1BWP7T $T=486520 672440 1 180 $X=475590 $Y=672205
X1307 36 265 6 5 19 DFQD1BWP7T $T=503880 695960 0 180 $X=492950 $Y=691750
X1308 102 331 6 5 237 DFQD1BWP7T $T=545320 711640 0 180 $X=534390 $Y=707430
X1309 102 412 6 5 292 DFQD1BWP7T $T=587320 719480 1 180 $X=576390 $Y=719245
X1310 102 402 6 5 300 DFQD1BWP7T $T=588440 711640 0 180 $X=577510 $Y=707430
X1311 102 338 6 5 374 DFQD1BWP7T $T=592360 735160 1 180 $X=581430 $Y=734925
X1312 102 429 6 5 423 DFQD1BWP7T $T=599640 703800 0 180 $X=588710 $Y=699590
X1313 102 316 6 5 8 DFQD1BWP7T $T=600760 711640 1 180 $X=589830 $Y=711405
X1314 102 432 6 5 15 DFQD1BWP7T $T=601320 688120 1 180 $X=590390 $Y=687885
X1315 102 433 6 5 290 DFQD1BWP7T $T=601880 656760 0 180 $X=590950 $Y=652550
X1316 102 436 6 5 72 DFQD1BWP7T $T=607480 680280 1 180 $X=596550 $Y=680045
X1317 102 448 6 5 93 DFQD1BWP7T $T=612520 664600 1 180 $X=601590 $Y=664365
X1318 51 50 6 5 47 190 197 MOAI22D0BWP7T $T=466920 617560 0 180 $X=462710 $Y=613350
X1319 51 73 6 5 210 193 47 MOAI22D0BWP7T $T=480920 633240 0 180 $X=476710 $Y=629030
X1320 51 111 6 5 47 349 389 MOAI22D0BWP7T $T=580600 601880 1 180 $X=576390 $Y=601645
X1321 51 119 6 5 333 416 47 MOAI22D0BWP7T $T=592360 617560 1 0 $X=592070 $Y=613350
X1322 276 341 350 351 358 6 5 XNR4D0BWP7T $T=534680 625400 0 0 $X=534390 $Y=625165
X1323 344 352 339 318 293 6 5 XNR4D0BWP7T $T=547560 672440 0 180 $X=534390 $Y=668230
X1324 359 307 344 343 317 6 5 XNR4D0BWP7T $T=547560 688120 0 180 $X=534390 $Y=683910
X1325 350 396 389 370 294 6 5 XNR4D0BWP7T $T=570520 601880 1 180 $X=557350 $Y=601645
X1326 257 230 293 65 301 6 5 XOR4D0BWP7T $T=503880 680280 1 0 $X=503590 $Y=676070
X1327 281 288 294 296 305 6 5 XOR4D0BWP7T $T=506120 617560 1 0 $X=505830 $Y=613350
X1328 291 250 318 319 287 6 5 XOR4D0BWP7T $T=515640 672440 1 0 $X=515350 $Y=668230
X1329 329 345 343 356 354 6 5 XOR4D0BWP7T $T=535800 735160 0 0 $X=535510 $Y=734925
X1330 104 348 370 373 334 6 5 XOR4D0BWP7T $T=546440 601880 1 0 $X=546150 $Y=597670
X1331 105 360 351 376 385 6 5 XOR4D0BWP7T $T=547560 625400 0 0 $X=547270 $Y=625165
X1332 72 6 5 69 CKND1BWP7T $T=479800 735160 1 180 $X=477830 $Y=734925
X1333 107 6 5 247 CKND1BWP7T $T=565480 727320 0 180 $X=563510 $Y=723110
X1334 130 6 5 109 CKND1BWP7T $T=612520 601880 1 180 $X=610550 $Y=601645
X1335 123 6 5 68 CKND1BWP7T $T=622600 617560 1 180 $X=620630 $Y=617325
X1336 423 18 6 5 BUFFD1P5BWP7T $T=593480 672440 1 180 $X=590390 $Y=672205
X1337 109 5 10 406 6 NR2D0BWP7T $T=568280 617560 0 0 $X=567990 $Y=617325
X1338 332 340 5 96 6 292 342 AOI22D1BWP7T $T=534680 719480 0 0 $X=534390 $Y=719245
X1339 332 398 5 96 6 374 336 AOI22D1BWP7T $T=568840 743000 0 180 $X=564630 $Y=738790
X1340 91 6 5 47 INVD3BWP7T $T=508920 601880 0 180 $X=505270 $Y=597670
X1341 302 6 5 277 CKBD1BWP7T $T=517320 719480 0 180 $X=514790 $Y=715270
X1342 375 6 5 371 CKBD1BWP7T $T=555400 617560 1 0 $X=555110 $Y=613350
X1343 410 6 5 404 CKBD1BWP7T $T=576680 633240 1 0 $X=576390 $Y=629030
X1344 380 6 5 246 CKBD1BWP7T $T=583400 688120 0 180 $X=580870 $Y=683910
X1345 151 6 5 553 CKBD1BWP7T $T=685320 664600 1 0 $X=685030 $Y=660390
X1346 478 139 5 6 139 476 143 MAOI22D0BWP7T $T=634920 633240 0 0 $X=634630 $Y=633005
X1347 530 159 5 6 159 535 457 MAOI22D0BWP7T $T=677480 641080 0 180 $X=673270 $Y=636870
X1348 567 159 5 6 159 576 456 MAOI22D0BWP7T $T=702680 648920 0 0 $X=702390 $Y=648685
X1349 555 159 5 6 159 550 324 MAOI22D0BWP7T $T=706600 703800 0 180 $X=702390 $Y=699590
X1350 577 159 5 6 159 593 440 MAOI22D0BWP7T $T=710520 656760 0 0 $X=710230 $Y=656525
X1351 599 159 5 6 159 609 405 MAOI22D0BWP7T $T=729560 688120 1 180 $X=725350 $Y=687885
X1352 611 159 5 6 159 615 323 MAOI22D0BWP7T $T=737960 719480 0 180 $X=733750 $Y=715270
X1353 603 139 5 6 173 617 169 MAOI22D0BWP7T $T=738520 609720 1 180 $X=734310 $Y=609485
X1354 612 139 5 6 173 618 162 MAOI22D0BWP7T $T=738520 617560 1 180 $X=734310 $Y=617325
X1355 608 159 5 6 159 619 431 MAOI22D0BWP7T $T=738520 672440 1 180 $X=734310 $Y=672205
X1356 613 159 5 6 159 616 413 MAOI22D0BWP7T $T=738520 735160 1 180 $X=734310 $Y=734925
X1357 274 328 276 5 6 357 OA21D0BWP7T $T=555400 648920 1 180 $X=551750 $Y=648685
X1358 60 369 359 5 6 311 OA21D0BWP7T $T=555960 727320 1 180 $X=552310 $Y=727085
X1359 325 314 8 332 96 5 6 AOI22D0BWP7T $T=525160 735160 1 0 $X=524870 $Y=730950
X1360 399 393 300 332 96 5 6 AOI22D0BWP7T $T=567720 711640 1 180 $X=564070 $Y=711405
X1361 106 392 332 325 401 5 6 AOI22D0BWP7T $T=565480 735160 0 0 $X=565190 $Y=734925
X1362 419 421 18 332 96 5 6 AOI22D0BWP7T $T=587880 695960 1 180 $X=584230 $Y=695725
X1363 426 425 15 332 96 5 6 AOI22D0BWP7T $T=592360 680280 1 180 $X=588710 $Y=680045
X1364 106 417 332 340 442 5 6 AOI22D0BWP7T $T=604120 719480 0 0 $X=603830 $Y=719245
X1365 444 443 72 332 96 5 6 AOI22D0BWP7T $T=609160 688120 1 180 $X=605510 $Y=687885
X1366 106 450 332 399 455 5 6 AOI22D0BWP7T $T=609160 711640 0 0 $X=608870 $Y=711405
X1367 462 460 93 332 96 5 6 AOI22D0BWP7T $T=622040 656760 0 180 $X=618390 $Y=652550
X1368 106 438 332 398 463 5 6 AOI22D0BWP7T $T=618680 727320 1 0 $X=618390 $Y=723110
X1369 135 464 332 442 467 5 6 AOI22D0BWP7T $T=623720 719480 1 0 $X=623430 $Y=715270
X1370 135 466 332 401 469 5 6 AOI22D0BWP7T $T=625960 727320 1 0 $X=625670 $Y=723110
X1371 106 465 332 462 471 5 6 AOI22D0BWP7T $T=627080 656760 1 0 $X=626790 $Y=652550
X1372 106 454 332 419 479 5 6 AOI22D0BWP7T $T=627080 695960 0 0 $X=626790 $Y=695725
X1373 135 473 332 455 475 5 6 AOI22D0BWP7T $T=631000 719480 1 0 $X=630710 $Y=715270
X1374 135 477 332 463 481 5 6 AOI22D0BWP7T $T=633800 727320 1 0 $X=633510 $Y=723110
X1375 135 483 332 471 482 5 6 AOI22D0BWP7T $T=642200 641080 1 180 $X=638550 $Y=640845
X1376 106 480 332 426 487 5 6 AOI22D0BWP7T $T=638840 680280 0 0 $X=638550 $Y=680045
X1377 106 472 332 444 490 5 6 AOI22D0BWP7T $T=639960 688120 1 0 $X=639670 $Y=683910
X1378 147 492 138 497 478 5 6 AOI22D0BWP7T $T=647800 617560 0 180 $X=644150 $Y=613350
X1379 135 498 332 487 503 5 6 AOI22D0BWP7T $T=646120 680280 1 0 $X=645830 $Y=676070
X1380 481 499 332 146 507 5 6 AOI22D0BWP7T $T=646680 727320 1 0 $X=646390 $Y=723110
X1381 135 500 332 479 502 5 6 AOI22D0BWP7T $T=647240 695960 0 0 $X=646950 $Y=695725
X1382 135 501 332 490 506 5 6 AOI22D0BWP7T $T=648360 688120 1 0 $X=648070 $Y=683910
X1383 482 489 332 146 509 5 6 AOI22D0BWP7T $T=649480 648920 0 0 $X=649190 $Y=648685
X1384 152 516 138 512 520 5 6 AOI22D0BWP7T $T=660680 617560 1 0 $X=660390 $Y=613350
X1385 467 515 332 146 521 5 6 AOI22D0BWP7T $T=660680 719480 0 0 $X=660390 $Y=719245
X1386 155 522 138 153 512 5 6 AOI22D0BWP7T $T=665720 601880 0 180 $X=662070 $Y=597670
X1387 150 513 332 509 528 5 6 AOI22D0BWP7T $T=662360 648920 1 0 $X=662070 $Y=644710
X1388 156 526 138 524 497 5 6 AOI22D0BWP7T $T=669080 617560 0 180 $X=665430 $Y=613350
X1389 154 525 332 528 530 5 6 AOI22D0BWP7T $T=666840 641080 1 0 $X=666550 $Y=636870
X1390 150 531 332 507 527 5 6 AOI22D0BWP7T $T=671320 719480 1 180 $X=667670 $Y=719245
X1391 158 532 138 520 524 5 6 AOI22D0BWP7T $T=673000 609720 1 180 $X=669350 $Y=609485
X1392 475 514 332 146 541 5 6 AOI22D0BWP7T $T=669640 703800 0 0 $X=669350 $Y=703565
X1393 502 518 332 146 539 5 6 AOI22D0BWP7T $T=673000 695960 1 0 $X=672710 $Y=691750
X1394 503 536 332 146 540 5 6 AOI22D0BWP7T $T=674120 664600 0 0 $X=673830 $Y=664365
X1395 506 537 332 146 544 5 6 AOI22D0BWP7T $T=678040 672440 0 0 $X=677750 $Y=672205
X1396 154 546 332 527 555 5 6 AOI22D0BWP7T $T=685320 719480 1 0 $X=685030 $Y=715270
X1397 469 554 332 146 558 5 6 AOI22D0BWP7T $T=686440 727320 0 0 $X=686150 $Y=727085
X1398 150 560 332 540 562 5 6 AOI22D0BWP7T $T=689800 680280 0 0 $X=689510 $Y=680045
X1399 154 561 332 562 567 5 6 AOI22D0BWP7T $T=692040 664600 1 0 $X=691750 $Y=660390
X1400 150 556 332 541 569 5 6 AOI22D0BWP7T $T=692600 711640 0 0 $X=692310 $Y=711405
X1401 152 552 138 165 573 5 6 AOI22D0BWP7T $T=693160 609720 0 0 $X=692870 $Y=609485
X1402 152 565 138 547 572 5 6 AOI22D0BWP7T $T=693160 617560 0 0 $X=692870 $Y=617325
X1403 150 568 332 544 571 5 6 AOI22D0BWP7T $T=693160 680280 1 0 $X=692870 $Y=676070
X1404 150 564 332 521 570 5 6 AOI22D0BWP7T $T=693160 727320 1 0 $X=692870 $Y=723110
X1405 155 559 138 161 547 5 6 AOI22D0BWP7T $T=702680 601880 1 0 $X=702390 $Y=597670
X1406 158 574 138 572 591 5 6 AOI22D0BWP7T $T=702680 625400 1 0 $X=702390 $Y=621190
X1407 154 575 332 571 577 5 6 AOI22D0BWP7T $T=702680 664600 1 0 $X=702390 $Y=660390
X1408 150 578 332 558 587 5 6 AOI22D0BWP7T $T=705480 719480 0 0 $X=705190 $Y=719245
X1409 158 588 138 573 592 5 6 AOI22D0BWP7T $T=710520 617560 0 0 $X=710230 $Y=617325
X1410 156 594 138 591 596 5 6 AOI22D0BWP7T $T=713320 625400 1 0 $X=713030 $Y=621190
X1411 150 585 332 539 597 5 6 AOI22D0BWP7T $T=713880 680280 0 0 $X=713590 $Y=680045
X1412 154 589 332 569 599 5 6 AOI22D0BWP7T $T=718360 688120 0 0 $X=718070 $Y=687885
X1413 154 598 332 587 611 5 6 AOI22D0BWP7T $T=719480 703800 0 0 $X=719190 $Y=703565
X1414 147 600 138 596 603 5 6 AOI22D0BWP7T $T=721160 617560 1 0 $X=720870 $Y=613350
X1415 156 601 138 592 607 5 6 AOI22D0BWP7T $T=722840 625400 1 0 $X=722550 $Y=621190
X1416 154 605 332 597 608 5 6 AOI22D0BWP7T $T=722840 680280 0 0 $X=722550 $Y=680045
X1417 154 610 332 570 613 5 6 AOI22D0BWP7T $T=726200 735160 0 0 $X=725910 $Y=734925
X1418 147 614 138 607 612 5 6 AOI22D0BWP7T $T=729000 617560 0 0 $X=728710 $Y=617325
X1419 6 5 ICV_41 $T=461320 633240 0 0 $X=461030 $Y=633005
X1420 6 5 ICV_41 $T=477000 633240 0 0 $X=476710 $Y=633005
X1421 6 5 ICV_41 $T=511720 695960 0 0 $X=511430 $Y=695725
X1422 6 5 ICV_41 $T=519560 641080 1 0 $X=519270 $Y=636870
X1423 6 5 ICV_41 $T=534120 719480 1 0 $X=533830 $Y=715270
X1424 6 5 ICV_41 $T=560440 625400 0 0 $X=560150 $Y=625165
X1425 6 5 ICV_41 $T=560440 672440 1 0 $X=560150 $Y=668230
X1426 6 5 ICV_41 $T=560440 688120 1 0 $X=560150 $Y=683910
X1427 6 5 ICV_41 $T=576120 656760 1 0 $X=575830 $Y=652550
X1428 6 5 ICV_41 $T=576120 664600 0 0 $X=575830 $Y=664365
X1429 6 5 ICV_41 $T=576120 688120 0 0 $X=575830 $Y=687885
X1430 6 5 ICV_41 $T=618120 625400 0 0 $X=617830 $Y=625165
X1431 6 5 ICV_41 $T=618120 680280 0 0 $X=617830 $Y=680045
X1432 6 5 ICV_41 $T=636040 656760 0 0 $X=635750 $Y=656525
X1433 6 5 ICV_41 $T=643880 656760 1 0 $X=643590 $Y=652550
X1434 6 5 ICV_41 $T=645560 641080 1 0 $X=645270 $Y=636870
X1435 6 5 ICV_41 $T=645560 727320 0 0 $X=645270 $Y=727085
X1436 6 5 ICV_41 $T=660120 648920 0 0 $X=659830 $Y=648685
X1437 6 5 ICV_41 $T=678040 617560 0 0 $X=677750 $Y=617325
X1438 6 5 ICV_41 $T=678040 711640 0 0 $X=677750 $Y=711405
X1439 6 5 ICV_41 $T=679160 727320 1 0 $X=678870 $Y=723110
X1440 6 5 ICV_41 $T=687560 672440 1 0 $X=687270 $Y=668230
X1441 6 5 ICV_41 $T=702120 743000 1 0 $X=701830 $Y=738790
X1442 6 5 ICV_41 $T=720040 656760 1 0 $X=719750 $Y=652550
X1443 6 5 ICV_41 $T=727880 648920 1 0 $X=727590 $Y=644710
X1444 6 5 ICV_41 $T=727880 695960 1 0 $X=727590 $Y=691750
X1445 6 5 ICV_41 $T=729000 727320 0 0 $X=728710 $Y=727085
X1446 6 5 ICV_41 $T=729560 656760 0 0 $X=729270 $Y=656525
X1447 6 5 ICV_37 $T=450120 601880 1 0 $X=449830 $Y=597670
X1448 6 5 ICV_37 $T=481480 617560 1 0 $X=481190 $Y=613350
X1449 6 5 ICV_37 $T=501080 688120 0 0 $X=500790 $Y=687885
X1450 6 5 ICV_37 $T=512840 695960 1 0 $X=512550 $Y=691750
X1451 6 5 ICV_37 $T=520680 743000 1 0 $X=520390 $Y=738790
X1452 6 5 ICV_37 $T=521800 735160 1 0 $X=521510 $Y=730950
X1453 6 5 ICV_37 $T=529640 672440 0 0 $X=529350 $Y=672205
X1454 6 5 ICV_37 $T=548680 735160 0 0 $X=548390 $Y=734925
X1455 6 5 ICV_37 $T=550360 695960 0 0 $X=550070 $Y=695725
X1456 6 5 ICV_37 $T=571640 695960 0 0 $X=571350 $Y=695725
X1457 6 5 ICV_37 $T=576120 672440 0 0 $X=575830 $Y=672205
X1458 6 5 ICV_37 $T=576120 688120 1 0 $X=575830 $Y=683910
X1459 6 5 ICV_37 $T=613640 719480 1 0 $X=613350 $Y=715270
X1460 6 5 ICV_37 $T=618120 680280 1 0 $X=617830 $Y=676070
X1461 6 5 ICV_37 $T=640520 617560 0 0 $X=640230 $Y=617325
X1462 6 5 ICV_37 $T=647800 633240 0 0 $X=647510 $Y=633005
X1463 6 5 ICV_37 $T=669080 680280 1 0 $X=668790 $Y=676070
X1464 6 5 ICV_37 $T=670200 641080 1 0 $X=669910 $Y=636870
X1465 6 5 ICV_37 $T=689240 695960 1 0 $X=688950 $Y=691750
X1466 6 5 ICV_37 $T=697640 680280 0 0 $X=697350 $Y=680045
X1467 6 5 ICV_37 $T=697640 719480 1 0 $X=697350 $Y=715270
X1468 6 5 ICV_37 $T=702120 672440 0 0 $X=701830 $Y=672205
X1469 6 5 ICV_37 $T=702120 719480 0 0 $X=701830 $Y=719245
X1470 6 5 ICV_37 $T=702120 727320 1 0 $X=701830 $Y=723110
X1471 6 5 ICV_37 $T=721720 688120 0 0 $X=721430 $Y=687885
X1472 6 5 ICV_37 $T=724520 695960 0 0 $X=724230 $Y=695725
X1473 6 5 ICV_37 $T=739640 664600 0 0 $X=739350 $Y=664365
X1474 6 5 ICV_43 $T=450120 680280 1 0 $X=449830 $Y=676070
X1475 6 5 ICV_43 $T=450120 743000 1 0 $X=449830 $Y=738790
X1476 6 5 ICV_43 $T=473080 656760 1 0 $X=472790 $Y=652550
X1477 6 5 ICV_43 $T=479800 735160 0 0 $X=479510 $Y=734925
X1478 6 5 ICV_43 $T=501080 625400 0 0 $X=500790 $Y=625165
X1479 6 5 ICV_43 $T=501080 680280 1 0 $X=500790 $Y=676070
X1480 6 5 ICV_43 $T=537480 601880 1 0 $X=537190 $Y=597670
X1481 6 5 ICV_43 $T=576120 672440 1 0 $X=575830 $Y=668230
X1482 6 5 ICV_43 $T=603000 672440 1 0 $X=602710 $Y=668230
X1483 6 5 ICV_43 $T=603000 680280 1 0 $X=602710 $Y=676070
X1484 6 5 ICV_43 $T=630440 656760 1 0 $X=630150 $Y=652550
X1485 6 5 ICV_43 $T=636040 648920 0 0 $X=635750 $Y=648685
X1486 6 5 ICV_43 $T=638280 703800 1 0 $X=637990 $Y=699590
X1487 6 5 ICV_43 $T=671320 664600 0 0 $X=671030 $Y=664365
X1488 6 5 ICV_43 $T=702120 648920 1 0 $X=701830 $Y=644710
X1489 6 5 ICV_43 $T=725080 727320 1 0 $X=724790 $Y=723110
X1490 6 5 ICV_52 $T=450120 735160 1 0 $X=449830 $Y=730950
X1491 6 5 ICV_52 $T=453480 735160 0 0 $X=453190 $Y=734925
X1492 6 5 ICV_52 $T=457960 695960 0 0 $X=457670 $Y=695725
X1493 6 5 ICV_52 $T=465800 727320 1 0 $X=465510 $Y=723110
X1494 6 5 ICV_52 $T=487080 719480 0 0 $X=486790 $Y=719245
X1495 6 5 ICV_52 $T=502760 641080 1 0 $X=502470 $Y=636870
X1496 6 5 ICV_52 $T=511720 672440 1 0 $X=511430 $Y=668230
X1497 6 5 ICV_52 $T=529080 719480 0 0 $X=528790 $Y=719245
X1498 6 5 ICV_52 $T=545320 727320 1 0 $X=545030 $Y=723110
X1499 6 5 ICV_52 $T=571080 641080 0 0 $X=570790 $Y=640845
X1500 6 5 ICV_52 $T=576120 680280 0 0 $X=575830 $Y=680045
X1501 6 5 ICV_52 $T=585080 703800 1 0 $X=584790 $Y=699590
X1502 6 5 ICV_52 $T=597960 641080 1 0 $X=597670 $Y=636870
X1503 6 5 ICV_52 $T=622040 727320 1 0 $X=621750 $Y=723110
X1504 6 5 ICV_52 $T=660120 641080 1 0 $X=659830 $Y=636870
X1505 6 5 ICV_52 $T=678040 719480 1 0 $X=677750 $Y=715270
X1506 108 5 10 391 6 NR2XD0BWP7T $T=567160 633240 0 0 $X=566870 $Y=633005
X1507 6 5 ICV_38 $T=486520 641080 1 0 $X=486230 $Y=636870
X1508 6 5 ICV_38 $T=486520 672440 0 0 $X=486230 $Y=672205
X1509 6 5 ICV_38 $T=486520 735160 1 0 $X=486230 $Y=730950
X1510 6 5 ICV_38 $T=528520 633240 1 0 $X=528230 $Y=629030
X1511 6 5 ICV_38 $T=528520 641080 0 0 $X=528230 $Y=640845
X1512 6 5 ICV_38 $T=528520 680280 0 0 $X=528230 $Y=680045
X1513 6 5 ICV_38 $T=528520 695960 0 0 $X=528230 $Y=695725
X1514 6 5 ICV_38 $T=528520 735160 1 0 $X=528230 $Y=730950
X1515 6 5 ICV_38 $T=528520 743000 1 0 $X=528230 $Y=738790
X1516 6 5 ICV_38 $T=570520 617560 0 0 $X=570230 $Y=617325
X1517 6 5 ICV_38 $T=570520 648920 0 0 $X=570230 $Y=648685
X1518 6 5 ICV_38 $T=570520 680280 0 0 $X=570230 $Y=680045
X1519 6 5 ICV_38 $T=570520 695960 1 0 $X=570230 $Y=691750
X1520 6 5 ICV_38 $T=570520 703800 1 0 $X=570230 $Y=699590
X1521 6 5 ICV_38 $T=570520 727320 1 0 $X=570230 $Y=723110
X1522 6 5 ICV_38 $T=612520 601880 0 0 $X=612230 $Y=601645
X1523 6 5 ICV_38 $T=612520 609720 1 0 $X=612230 $Y=605510
X1524 6 5 ICV_38 $T=612520 641080 1 0 $X=612230 $Y=636870
X1525 6 5 ICV_38 $T=612520 695960 0 0 $X=612230 $Y=695725
X1526 6 5 ICV_38 $T=612520 711640 0 0 $X=612230 $Y=711405
X1527 6 5 ICV_38 $T=612520 735160 1 0 $X=612230 $Y=730950
X1528 6 5 ICV_38 $T=654520 633240 0 0 $X=654230 $Y=633005
X1529 6 5 ICV_38 $T=654520 641080 0 0 $X=654230 $Y=640845
X1530 6 5 ICV_38 $T=654520 703800 0 0 $X=654230 $Y=703565
X1531 6 5 ICV_38 $T=696520 695960 1 0 $X=696230 $Y=691750
X1532 6 5 ICV_38 $T=696520 727320 1 0 $X=696230 $Y=723110
X1533 6 5 ICV_45 $T=450120 641080 1 0 $X=449830 $Y=636870
X1534 6 5 ICV_45 $T=455720 735160 1 0 $X=455430 $Y=730950
X1535 6 5 ICV_45 $T=463560 609720 0 0 $X=463270 $Y=609485
X1536 6 5 ICV_45 $T=463560 680280 1 0 $X=463270 $Y=676070
X1537 6 5 ICV_45 $T=464120 601880 1 0 $X=463830 $Y=597670
X1538 6 5 ICV_45 $T=502760 672440 0 0 $X=502470 $Y=672205
X1539 6 5 ICV_45 $T=534120 617560 0 0 $X=533830 $Y=617325
X1540 6 5 ICV_45 $T=534120 703800 1 0 $X=533830 $Y=699590
X1541 6 5 ICV_45 $T=576120 680280 1 0 $X=575830 $Y=676070
X1542 6 5 ICV_45 $T=583400 688120 1 0 $X=583110 $Y=683910
X1543 6 5 ICV_45 $T=588440 711640 1 0 $X=588150 $Y=707430
X1544 6 5 ICV_45 $T=589560 609720 0 0 $X=589270 $Y=609485
X1545 6 5 ICV_45 $T=618120 703800 0 0 $X=617830 $Y=703565
X1546 6 5 ICV_45 $T=660120 633240 0 0 $X=659830 $Y=633005
X1547 6 5 ICV_45 $T=660120 688120 0 0 $X=659830 $Y=687885
X1548 6 5 ICV_45 $T=671880 625400 1 0 $X=671590 $Y=621190
X1549 6 5 ICV_45 $T=708840 664600 1 0 $X=708550 $Y=660390
X1550 6 5 ICV_45 $T=712760 664600 0 0 $X=712470 $Y=664365
X1551 6 5 ICV_45 $T=715000 688120 1 0 $X=714710 $Y=683910
X1552 124 6 5 120 BUFFD3BWP7T $T=597400 727320 0 180 $X=593190 $Y=723110
X1553 172 6 5 171 BUFFD3BWP7T $T=723400 719480 0 180 $X=719190 $Y=715270
X1554 622 6 5 170 BUFFD3BWP7T $T=737960 656760 0 180 $X=733750 $Y=652550
X1555 277 372 6 5 346 362 IAO21D0BWP7T $T=567160 695960 0 180 $X=563510 $Y=691750
X1556 290 390 6 5 386 388 IAO21D0BWP7T $T=582280 672440 0 180 $X=578630 $Y=668230
X1557 85 371 262 5 6 377 AN3D1BWP7T $T=553160 656760 0 0 $X=552870 $Y=656525
X1558 85 404 277 5 6 346 AN3D1BWP7T $T=570520 695960 0 180 $X=566870 $Y=691750
X1559 85 384 290 5 6 386 AN3D1BWP7T $T=580040 680280 0 0 $X=579750 $Y=680045
X1560 144 130 434 5 6 129 AN3D1BWP7T $T=638840 601880 1 180 $X=635190 $Y=601645
X1561 157 5 102 6 CKND12BWP7T $T=669640 672440 0 180 $X=660390 $Y=668230
X1562 36 225 60 6 5 DFQD2BWP7T $T=483720 664600 0 180 $X=472230 $Y=660390
X1563 136 6 5 332 BUFFD5BWP7T $T=627080 641080 0 0 $X=626790 $Y=640845
X1564 136 6 5 138 BUFFD5BWP7T $T=627640 617560 1 0 $X=627350 $Y=613350
X1565 171 323 553 6 5 ND2D2BWP7T $T=692600 695960 1 0 $X=692310 $Y=691750
X1566 160 413 151 6 5 ND2D1P5BWP7T $T=678600 648920 1 180 $X=674390 $Y=648685
X1567 164 324 151 6 5 ND2D1P5BWP7T $T=687560 633240 0 0 $X=687270 $Y=633005
X1568 51 262 6 243 191 47 5 MOAI22D1BWP7T $T=497720 641080 1 180 $X=492950 $Y=640845
X1569 51 277 6 47 198 270 5 MOAI22D1BWP7T $T=506120 656760 0 180 $X=501350 $Y=652550
X1570 51 305 6 47 234 339 5 MOAI22D1BWP7T $T=539160 656760 0 180 $X=534390 $Y=652550
X1571 51 434 6 47 430 428 5 MOAI22D1BWP7T $T=606360 641080 1 180 $X=601590 $Y=640845
X1572 51 148 6 47 439 452 5 MOAI22D1BWP7T $T=652840 601880 0 180 $X=648070 $Y=597670
X1573 262 381 5 377 322 6 IAO21D1BWP7T $T=556520 656760 0 0 $X=556230 $Y=656525
X1574 434 449 5 129 127 6 IAO21D1BWP7T $T=610840 601880 1 180 $X=606630 $Y=601645
X1575 323 96 5 314 316 6 OAI21D1BWP7T $T=524600 719480 1 180 $X=520950 $Y=719245
X1576 324 96 5 336 338 6 OAI21D1BWP7T $T=525160 727320 1 0 $X=524870 $Y=723110
X1577 106 323 5 392 394 6 OAI21D1BWP7T $T=565480 727320 0 0 $X=565190 $Y=727085
X1614 6 5 ICV_51 $T=489320 625400 1 0 $X=489030 $Y=621190
X1615 6 5 ICV_51 $T=489320 688120 0 0 $X=489030 $Y=687885
X1616 6 5 ICV_51 $T=489320 703800 1 0 $X=489030 $Y=699590
X1617 6 5 ICV_51 $T=531320 633240 0 0 $X=531030 $Y=633005
X1618 6 5 ICV_51 $T=531320 695960 1 0 $X=531030 $Y=691750
X1619 6 5 ICV_51 $T=573320 727320 0 0 $X=573030 $Y=727085
X1620 6 5 ICV_51 $T=573320 743000 1 0 $X=573030 $Y=738790
X1621 6 5 ICV_51 $T=615320 680280 1 0 $X=615030 $Y=676070
X1622 6 5 ICV_51 $T=615320 711640 1 0 $X=615030 $Y=707430
X1623 6 5 ICV_51 $T=615320 735160 0 0 $X=615030 $Y=734925
X1624 6 5 ICV_51 $T=657320 601880 1 0 $X=657030 $Y=597670
X1625 6 5 ICV_51 $T=657320 648920 1 0 $X=657030 $Y=644710
X1626 6 5 ICV_51 $T=657320 648920 0 0 $X=657030 $Y=648685
X1627 6 5 ICV_51 $T=657320 656760 1 0 $X=657030 $Y=652550
X1628 6 5 ICV_51 $T=657320 703800 1 0 $X=657030 $Y=699590
X1629 6 5 ICV_51 $T=657320 719480 1 0 $X=657030 $Y=715270
X1630 6 5 ICV_51 $T=699320 641080 1 0 $X=699030 $Y=636870
X1631 6 5 ICV_51 $T=699320 656760 1 0 $X=699030 $Y=652550
X1632 6 5 ICV_51 $T=699320 695960 0 0 $X=699030 $Y=695725
X1633 6 5 ICV_51 $T=699320 719480 0 0 $X=699030 $Y=719245
X1634 6 5 ICV_39 $T=486520 617560 1 0 $X=486230 $Y=613350
X1635 6 5 ICV_39 $T=486520 641080 0 0 $X=486230 $Y=640845
X1636 6 5 ICV_39 $T=738520 601880 0 0 $X=738230 $Y=601645
X1637 6 5 ICV_39 $T=738520 609720 0 0 $X=738230 $Y=609485
X1638 6 5 ICV_39 $T=738520 617560 0 0 $X=738230 $Y=617325
X1639 6 5 ICV_39 $T=738520 625400 1 0 $X=738230 $Y=621190
X1640 6 5 ICV_39 $T=738520 633240 1 0 $X=738230 $Y=629030
X1641 6 5 ICV_39 $T=738520 641080 0 0 $X=738230 $Y=640845
X1642 6 5 ICV_39 $T=738520 672440 1 0 $X=738230 $Y=668230
X1643 6 5 ICV_39 $T=738520 672440 0 0 $X=738230 $Y=672205
X1644 6 5 ICV_39 $T=738520 680280 0 0 $X=738230 $Y=680045
X1645 6 5 ICV_39 $T=738520 688120 0 0 $X=738230 $Y=687885
X1646 6 5 ICV_39 $T=738520 695960 0 0 $X=738230 $Y=695725
X1647 6 5 ICV_39 $T=738520 711640 1 0 $X=738230 $Y=707430
X1648 6 5 ICV_39 $T=738520 727320 1 0 $X=738230 $Y=723110
X1649 6 5 ICV_39 $T=738520 735160 0 0 $X=738230 $Y=734925
X1650 6 5 ICV_42 $T=450120 609720 1 0 $X=449830 $Y=605510
X1651 6 5 ICV_42 $T=492120 735160 1 0 $X=491830 $Y=730950
X1652 6 5 ICV_42 $T=515640 633240 0 0 $X=515350 $Y=633005
X1653 6 5 ICV_42 $T=516760 625400 0 0 $X=516470 $Y=625165
X1654 6 5 ICV_42 $T=516760 680280 1 0 $X=516470 $Y=676070
X1655 6 5 ICV_42 $T=517320 719480 1 0 $X=517030 $Y=715270
X1656 6 5 ICV_42 $T=539160 656760 1 0 $X=538870 $Y=652550
X1657 6 5 ICV_42 $T=559320 601880 1 0 $X=559030 $Y=597670
X1658 6 5 ICV_42 $T=576120 609720 1 0 $X=575830 $Y=605510
X1659 6 5 ICV_42 $T=576120 617560 1 0 $X=575830 $Y=613350
X1660 6 5 ICV_42 $T=576120 617560 0 0 $X=575830 $Y=617325
X1661 6 5 ICV_42 $T=576120 727320 1 0 $X=575830 $Y=723110
X1662 6 5 ICV_42 $T=587320 719480 0 0 $X=587030 $Y=719245
X1663 6 5 ICV_42 $T=599640 703800 1 0 $X=599350 $Y=699590
X1664 6 5 ICV_42 $T=618120 672440 1 0 $X=617830 $Y=668230
X1665 6 5 ICV_42 $T=702120 719480 1 0 $X=701830 $Y=715270
X1666 6 5 ICV_42 $T=702120 727320 0 0 $X=701830 $Y=727085
X1667 6 5 ICV_42 $T=725640 625400 0 0 $X=725350 $Y=625165
X1668 6 5 ICV_42 $T=726760 719480 0 0 $X=726470 $Y=719245
X1669 6 5 ICV_42 $T=727320 609720 1 0 $X=727030 $Y=605510
X1670 6 5 ICV_42 $T=727320 711640 0 0 $X=727030 $Y=711405
X1671 237 6 5 26 CKND0BWP7T $T=454600 743000 0 180 $X=452630 $Y=738790
X1672 6 5 ICV_48 $T=450120 672440 0 0 $X=449830 $Y=672205
X1673 6 5 ICV_48 $T=492120 617560 0 0 $X=491830 $Y=617325
X1674 6 5 ICV_48 $T=507240 735160 0 0 $X=506950 $Y=734925
X1675 6 5 ICV_48 $T=508360 648920 0 0 $X=508070 $Y=648685
X1676 6 5 ICV_48 $T=534120 633240 1 0 $X=533830 $Y=629030
X1677 6 5 ICV_48 $T=576120 703800 0 0 $X=575830 $Y=703565
X1678 6 5 ICV_48 $T=576120 719480 1 0 $X=575830 $Y=715270
X1679 6 5 ICV_48 $T=576120 735160 1 0 $X=575830 $Y=730950
X1680 6 5 ICV_48 $T=618120 664600 1 0 $X=617830 $Y=660390
X1681 6 5 ICV_48 $T=633240 688120 0 0 $X=632950 $Y=687885
X1682 6 5 ICV_48 $T=660120 664600 1 0 $X=659830 $Y=660390
X1683 6 5 ICV_48 $T=660120 727320 0 0 $X=659830 $Y=727085
X1684 6 5 ICV_48 $T=663480 609720 1 0 $X=663190 $Y=605510
X1685 6 5 ICV_48 $T=702120 601880 0 0 $X=701830 $Y=601645
X1686 6 5 ICV_48 $T=702120 633240 1 0 $X=701830 $Y=629030
X1687 6 5 ICV_48 $T=702120 641080 0 0 $X=701830 $Y=640845
.ENDS
***************************************
.SUBCKT __$$VIA34_520_520_60_21
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_72 2 3 4 5 6 7 9 10 11 12 13
** N=14 EP=11 IP=154 FDC=490
*.SEEDPROM
X52 6 2 7 7 3 10 11 11 10 9 10 7 PDDW0208CDG $T=530170 0 0 0 $X=529570 $Y=0
X53 6 2 7 7 4 10 11 11 10 12 10 7 PDDW0208CDG $T=610200 0 0 0 $X=609600 $Y=0
X54 6 2 7 7 5 10 11 11 10 13 10 7 PDDW0208CDG $T=690240 0 0 0 $X=689640 $Y=0
X55 6 2 7 7 7 PVDD1CDG $T=450135 0 0 0 $X=449535 $Y=0
.ENDS
***************************************
.SUBCKT ICV_34 2 3 4 5 6 7 8 10 11 12 14
** N=27 EP=11 IP=184 FDC=490
*.SEEDPROM
M0 6 17 16 6 PD L=1.6e-06 W=7.5e-07 $X=702380 $Y=810110 $D=17
M1 7 23 27 6 PD L=6e-07 W=5e-06 $X=710220 $Y=812390 $D=17
M2 23 16 27 6 PD L=6e-07 W=4.5e-06 $X=714690 $Y=812890 $D=17
M3 27 16 23 6 PD L=6e-07 W=4.5e-06 $X=716290 $Y=812890 $D=17
M4 23 22 6 6 PD L=6e-07 W=1.5e-06 $X=717890 $Y=809890 $D=17
M5 6 16 27 6 PD L=6e-07 W=4.5e-06 $X=717890 $Y=812890 $D=17
M6 6 22 23 6 PD L=6e-07 W=1.5e-06 $X=719490 $Y=809890 $D=17
M7 27 16 6 6 PD L=6e-07 W=4.5e-06 $X=719490 $Y=812890 $D=17
X44 6 7 18 19 20 21 5 7 HBK183_POSTDRV_PDUW0208SCDG_S $T=770240 900000 0 180 $X=689640 $Y=807690
X45 6 2 7 11 18 19 10 20 21 10 11 22 14 24 23 11 17 16 5 7 HBK183_PREDRV $T=770240 818990 0 180 $X=689640 $Y=780000
X51 7 22 6 23 16 HBK183_SCH_CELL $T=722190 818410 0 180 $X=707400 $Y=791530
X54 6 2 7 7 3 10 8 11 10 25 10 7 PDDW0208CDG $T=610170 900000 0 180 $X=529570 $Y=780000
X55 6 2 7 7 4 10 12 11 10 26 10 7 PDDW0208CDG $T=690200 900000 0 180 $X=609600 $Y=780000
X69 6 2 7 7 7 PVDD1CDG $T=530135 900000 0 180 $X=449535 $Y=780000
.ENDS
***************************************
.SUBCKT ICV_26 1 2 3 4 5 6 7
** N=8 EP=7 IP=13 FDC=145
*.SEEDPROM
X0 1 2 3 3 7 4 5 5 4 6 4 3 PDDW0208CDG $T=0 0 0 0 $X=-600 $Y=0
.ENDS
***************************************
.SUBCKT ICV_24 1 2 3 4 5 6 7
** N=8 EP=7 IP=13 FDC=145
*.SEEDPROM
X0 1 2 3 3 7 4 5 5 4 6 4 3 PDDW0208CDG $T=0 0 0 0 $X=-600 $Y=0
.ENDS
***************************************
.SUBCKT ICV_22 1 3
** N=4 EP=2 IP=6 FDC=60
*.SEEDPROM
X0 1 3 3 3 PVDD2CDG $T=0 0 0 0 $X=-600 $Y=0
.ENDS
***************************************
.SUBCKT ICV_17 1 2 3
** N=4 EP=3 IP=6 FDC=55
*.SEEDPROM
X0 1 2 3 3 3 PVDD1CDG $T=0 0 0 0 $X=-600 $Y=0
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4 5 6 7
** N=8 EP=7 IP=13 FDC=145
*.SEEDPROM
X0 1 2 3 3 7 5 6 6 5 4 5 3 PDDW0208CDG $T=0 0 0 0 $X=-600 $Y=0
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6 7
** N=8 EP=7 IP=13 FDC=145
*.SEEDPROM
X0 1 2 3 3 7 4 6 6 4 5 4 3 PDDW0208CDG $T=0 0 0 0 $X=-600 $Y=0
.ENDS
***************************************
.SUBCKT systolic_array p_shift_out<3> VDD p_shift_out<0> p_shift_in<4> p_shift_in<3> clk_p en_p VDDPST VSS p_shift_out<4> p_shift_out<2> p_shift_out<1> p_shift_out<5> p_shift_out<6> p_shift_in<2> p_shift_in<1> p_shift_in<0> p_shift_in<7> p_shift_in<6> p_shift_in<5>
+ p_shift_out<7> ack_p rstn_p
** N=987 EP=23 IP=2284 FDC=113190
D0 VSS VDDPST pnwdio_5_iso AREA=4.37643e-08 pj=0.0135966 $X=36190 $Y=124715 $D=112
D1 VSS VDD pnwdio_iso AREA=1.27584e-08 pj=0.00564005 $X=110050 $Y=128725 $D=114
D2 VSS VDD pnwdio_iso AREA=2.53754e-09 pj=0.00119151 $X=154710 $Y=235175 $D=114
D3 VSS VDD pnwdio_iso AREA=2.54139e-09 pj=0.00119148 $X=154710 $Y=352775 $D=114
D4 VSS VDD pnwdio_iso AREA=2.53698e-09 pj=0.00119121 $X=154710 $Y=478215 $D=114
D5 VSS VDD pnwdio_iso AREA=2.53528e-09 pj=0.00119076 $X=154710 $Y=595815 $D=114
D6 VSS VDD pnwdio_iso AREA=2.53661e-09 pj=0.00119184 $X=154710 $Y=156775 $D=114
D7 VSS VDD pnwdio_iso AREA=2.5355e-09 pj=0.00119094 $X=154710 $Y=172455 $D=114
D8 VSS VDD pnwdio_iso AREA=2.53565e-09 pj=0.00119106 $X=154710 $Y=188135 $D=114
D9 VSS VDD pnwdio_iso AREA=2.53558e-09 pj=0.001191 $X=154710 $Y=195975 $D=114
D10 VSS VDD pnwdio_iso AREA=2.53535e-09 pj=0.00119082 $X=154710 $Y=203815 $D=114
D11 VSS VDD pnwdio_iso AREA=2.5358e-09 pj=0.00119118 $X=154710 $Y=211655 $D=114
D12 VSS VDD pnwdio_iso AREA=2.53491e-09 pj=0.00119046 $X=154710 $Y=219495 $D=114
D13 VSS VDD pnwdio_iso AREA=2.53788e-09 pj=0.00119187 $X=154710 $Y=227335 $D=114
D14 VSS VDD pnwdio_iso AREA=2.53499e-09 pj=0.00119052 $X=154710 $Y=164615 $D=114
D15 VSS VDD pnwdio_iso AREA=2.53528e-09 pj=0.00119076 $X=154710 $Y=180295 $D=114
D16 VSS VDD pnwdio_iso AREA=2.53565e-09 pj=0.00119106 $X=154710 $Y=243015 $D=114
D17 VSS VDD pnwdio_iso AREA=2.53587e-09 pj=0.00119124 $X=154710 $Y=250855 $D=114
D18 VSS VDD pnwdio_iso AREA=2.53883e-09 pj=0.00119178 $X=154710 $Y=258695 $D=114
D19 VSS VDD pnwdio_iso AREA=2.5358e-09 pj=0.00119118 $X=154710 $Y=266535 $D=114
D20 VSS VDD pnwdio_iso AREA=2.5355e-09 pj=0.00119094 $X=154710 $Y=274375 $D=114
D21 VSS VDD pnwdio_iso AREA=2.53558e-09 pj=0.001191 $X=154710 $Y=282215 $D=114
D22 VSS VDD pnwdio_iso AREA=2.53543e-09 pj=0.00119088 $X=154710 $Y=290055 $D=114
D23 VSS VDD pnwdio_iso AREA=2.53587e-09 pj=0.00119124 $X=154710 $Y=297895 $D=114
D24 VSS VDD pnwdio_iso AREA=2.53528e-09 pj=0.00119076 $X=154710 $Y=305735 $D=114
D25 VSS VDD pnwdio_iso AREA=2.53706e-09 pj=0.00119127 $X=154710 $Y=313575 $D=114
D26 VSS VDD pnwdio_iso AREA=2.53521e-09 pj=0.0011907 $X=154710 $Y=321415 $D=114
D27 VSS VDD pnwdio_iso AREA=2.53728e-09 pj=0.00119145 $X=154710 $Y=329255 $D=114
D28 VSS VDD pnwdio_iso AREA=2.53528e-09 pj=0.00119076 $X=154710 $Y=337095 $D=114
D29 VSS VDD pnwdio_iso AREA=2.53958e-09 pj=0.00119162 $X=154710 $Y=344935 $D=114
D30 VSS VDD pnwdio_iso AREA=2.5355e-09 pj=0.00119094 $X=154710 $Y=360615 $D=114
D31 VSS VDD pnwdio_iso AREA=2.53535e-09 pj=0.00119082 $X=154710 $Y=368455 $D=114
D32 VSS VDD pnwdio_iso AREA=2.53565e-09 pj=0.00119106 $X=154710 $Y=376295 $D=114
D33 VSS VDD pnwdio_iso AREA=2.53544e-09 pj=0.00119161 $X=154710 $Y=384135 $D=114
D34 VSS VDD pnwdio_iso AREA=2.53796e-09 pj=0.00119165 $X=154710 $Y=391975 $D=114
D35 VSS VDD pnwdio_iso AREA=2.5383e-09 pj=0.00119156 $X=154710 $Y=399815 $D=114
D36 VSS VDD pnwdio_iso AREA=2.535e-09 pj=0.00119125 $X=154710 $Y=407655 $D=114
D37 VSS VDD pnwdio_iso AREA=2.53513e-09 pj=0.00119064 $X=154710 $Y=415495 $D=114
D38 VSS VDD pnwdio_iso AREA=2.53507e-09 pj=0.00119131 $X=154710 $Y=423335 $D=114
D39 VSS VDD pnwdio_iso AREA=2.54092e-09 pj=0.0011915 $X=154710 $Y=431175 $D=114
D40 VSS VDD pnwdio_iso AREA=2.53929e-09 pj=0.00119138 $X=154710 $Y=439015 $D=114
D41 VSS VDD pnwdio_iso AREA=2.53951e-09 pj=0.00119144 $X=154710 $Y=446855 $D=114
D42 VSS VDD pnwdio_iso AREA=2.53521e-09 pj=0.0011907 $X=154710 $Y=454695 $D=114
D43 VSS VDD pnwdio_iso AREA=2.53521e-09 pj=0.0011907 $X=154710 $Y=462535 $D=114
D44 VSS VDD pnwdio_iso AREA=2.53521e-09 pj=0.0011907 $X=154710 $Y=470375 $D=114
D45 VSS VDD pnwdio_iso AREA=2.53506e-09 pj=0.00119058 $X=154710 $Y=486055 $D=114
D46 VSS VDD pnwdio_iso AREA=2.53968e-09 pj=0.00119124 $X=154710 $Y=493895 $D=114
D47 VSS VDD pnwdio_iso AREA=2.53506e-09 pj=0.00119058 $X=154710 $Y=501735 $D=114
D48 VSS VDD pnwdio_iso AREA=2.53513e-09 pj=0.00119064 $X=154710 $Y=509575 $D=114
D49 VSS VDD pnwdio_iso AREA=2.53558e-09 pj=0.001191 $X=154710 $Y=517415 $D=114
D50 VSS VDD pnwdio_iso AREA=2.53572e-09 pj=0.00119112 $X=154710 $Y=525255 $D=114
D51 VSS VDD pnwdio_iso AREA=2.53558e-09 pj=0.001191 $X=154710 $Y=533095 $D=114
D52 VSS VDD pnwdio_iso AREA=2.53543e-09 pj=0.00119088 $X=154710 $Y=540935 $D=114
D53 VSS VDD pnwdio_iso AREA=2.53513e-09 pj=0.00119064 $X=154710 $Y=548775 $D=114
D54 VSS VDD pnwdio_iso AREA=2.53858e-09 pj=0.00119141 $X=154710 $Y=556615 $D=114
D55 VSS VDD pnwdio_iso AREA=2.53528e-09 pj=0.00119076 $X=154710 $Y=564455 $D=114
D56 VSS VDD pnwdio_iso AREA=2.53521e-09 pj=0.0011907 $X=154710 $Y=572295 $D=114
D57 VSS VDD pnwdio_iso AREA=2.53521e-09 pj=0.0011907 $X=154710 $Y=580135 $D=114
D58 VSS VDD pnwdio_iso AREA=2.53837e-09 pj=0.00119162 $X=154710 $Y=587975 $D=114
D59 VSS VDD pnwdio_iso AREA=2.53865e-09 pj=0.00119147 $X=154710 $Y=603655 $D=114
D60 VSS VDD pnwdio_iso AREA=2.53535e-09 pj=0.00119082 $X=154710 $Y=611495 $D=114
D61 VSS VDD pnwdio_iso AREA=2.53543e-09 pj=0.00119088 $X=154710 $Y=619335 $D=114
D62 VSS VDD pnwdio_iso AREA=2.53558e-09 pj=0.001191 $X=154710 $Y=627175 $D=114
D63 VSS VDD pnwdio_iso AREA=2.53543e-09 pj=0.00119088 $X=154710 $Y=635015 $D=114
D64 VSS VDD pnwdio_iso AREA=2.53543e-09 pj=0.00119088 $X=154710 $Y=642855 $D=114
D65 VSS VDD pnwdio_iso AREA=2.53737e-09 pj=0.00119145 $X=154710 $Y=650695 $D=114
D66 VSS VDD pnwdio_iso AREA=2.53513e-09 pj=0.00119064 $X=154710 $Y=658535 $D=114
D67 VSS VDD pnwdio_iso AREA=2.5372e-09 pj=0.00119139 $X=154710 $Y=666375 $D=114
D68 VSS VDD pnwdio_iso AREA=2.53513e-09 pj=0.00119064 $X=154710 $Y=674215 $D=114
D69 VSS VDD pnwdio_iso AREA=2.53543e-09 pj=0.00119088 $X=154710 $Y=682055 $D=114
D70 VSS VDD pnwdio_iso AREA=2.53558e-09 pj=0.001191 $X=154710 $Y=689895 $D=114
D71 VSS VDD pnwdio_iso AREA=2.53499e-09 pj=0.00119052 $X=154710 $Y=697735 $D=114
D72 VSS VDD pnwdio_iso AREA=2.53572e-09 pj=0.00119112 $X=154710 $Y=705575 $D=114
D73 VSS VDD pnwdio_iso AREA=2.53469e-09 pj=0.00119028 $X=154710 $Y=713415 $D=114
D74 VSS VDD pnwdio_iso AREA=2.53521e-09 pj=0.0011907 $X=154710 $Y=721255 $D=114
D75 VSS VDD pnwdio_iso AREA=2.53477e-09 pj=0.00119034 $X=154710 $Y=729095 $D=114
D76 VSS VDD pnwdio_iso AREA=2.53572e-09 pj=0.00119112 $X=154710 $Y=736935 $D=114
X83 clk_p en_p VDDPST VSS VDD 39 25 26 867 ICV_85 $T=0 0 0 0 $X=-25000 $Y=-25000
X88 VSS VDD 48 49 42 46 83 868 67 43 45 44 51 870 54 50 869 47 63 52
+ 872 867 877 57 77 53 55 64 56 60 59 871 58 61 62 163 93 876 75 65
+ 874 69 72 68 70 71 873 73 81 74 66 76 84 78 79 88 80 82 86 85
+ 97 91 87 90 92 714 96 89 98 99 101 100 875 94 95 103 105 113 106 123
+ 107 120 443 435 102 108 118 109 104 110 111 114 721 439 440 112 115 718 121 117
+ 127 116 125 726 436 712 122 119 723 724 733 717 128 124 727 878 126 716 713 728
+ 725 722 28 720 719 715
+ ICV_84 $T=0 0 0 0 $X=-25000 $Y=141500
X89 VSS VDD 872 139 135 130 881 868 46 131 42 132 136 883 138 133 134 147 880 879
+ 45 146 137 160 141 882 140 49 47 156 145 43 64 50 56 152 51 142 148 71
+ 52 53 54 163 55 870 144 57 59 150 871 155 62 63 149 60 58 143 151 158
+ 68 44 76 159 66 889 169 887 79 157 69 67 61 884 74 72 73 162 166 154
+ 153 164 75 48 165 167 77 70 161 87 168 885 80 170 203 172 177 171 179 184
+ 886 176 265 82 83 78 65 174 175 84 85 86 199 178 173 88 89 869 192 90
+ 186 182 183 91 93 180 98 202 733 94 99 215 95 200 103 114 191 185 96 81
+ 187 714 97 92 873 206 189 742 874 188 190 875 876 102 193 100 101 194 201 111
+ 104 195 196 750 197 106 198 888 877 209 109 207 110 213 108 105 204 112 205 113
+ 181 211 890 115 118 208 107 732 116 222 210 729 121 117 891 119 736 741 748 122
+ 738 217 212 214 218 125 220 123 219 221 216 124 878 126 745 223 749 420 740 225
+ 730 224 120 744 504 743 746 226 421 128 734 127 737 544 494 735 739 29 424 731
+ 747 30
+ ICV_83 $T=0 0 0 0 $X=-25000 $Y=241000
X90 VDD VSS VDDPST 872 130 227 879 893 46 230 240 228 892 133 229 232 134 880 132 234
+ 233 237 235 231 136 138 151 236 881 135 239 131 899 238 241 896 137 139 56 64
+ 882 883 163 242 243 141 153 244 142 143 907 245 144 146 145 140 246 147 164 902
+ 249 148 904 149 248 150 897 152 900 59 256 168 908 898 895 167 901 154 155 903
+ 157 250 894 156 158 906 159 160 253 252 161 165 905 254 162 247 258 255 271 269
+ 169 166 257 174 909 264 270 272 170 910 277 171 178 911 205 266 176 172 259 263
+ 175 173 265 886 261 260 180 177 273 885 262 267 268 251 179 181 185 184 182 192
+ 742 778 274 912 215 183 884 187 191 189 188 275 186 276 194 887 209 913 190 888
+ 204 196 279 197 195 281 284 283 278 914 280 286 774 291 282 287 915 199 388 285
+ 193 206 200 288 889 201 311 295 289 202 290 203 300 292 297 208 296 293 299 777
+ 766 781 207 890 294 575 298 307 212 770 302 771 210 303 213 768 214 222 316 304
+ 305 760 306 198 310 757 761 301 217 211 216 754 803 308 218 219 220 783 775 763
+ 776 779 312 224 313 916 320 562 221 315 753 223 32 314 767 317 765 784 782 769
+ 31 758 755 751 756 772 225 891 226 762 752 780 496 773 495 764 321 759
+ ICV_82 $T=0 0 0 0 $X=-25000 $Y=358600
X91 VDD VSS 893 250 247 902 325 892 324 228 233 327 230 323 919 227 918 330 326 231
+ 917 331 234 322 129 232 921 235 894 328 229 349 237 238 240 239 895 332 909 236
+ 905 333 345 336 351 341 922 241 334 243 896 897 335 337 901 903 353 924 244 329
+ 338 265 906 245 246 339 242 176 248 252 344 340 249 346 350 172 927 923 343 928
+ 253 361 926 260 920 352 925 251 355 258 347 342 254 358 256 360 257 261 259 255
+ 363 262 364 362 263 267 366 264 370 365 911 280 367 931 733 910 356 354 368 348
+ 268 275 929 371 930 908 169 269 375 359 357 270 912 376 377 276 373 932 369 378
+ 388 271 282 914 379 913 266 273 383 279 372 274 272 381 382 384 389 277 391 278
+ 394 380 398 385 397 281 790 386 933 402 287 935 934 285 387 284 399 936 798 939
+ 374 916 289 286 403 288 290 390 393 291 396 307 392 283 295 294 915 794 296 293
+ 299 297 300 303 292 400 395 301 401 938 298 937 405 304 789 404 803 305 788 306
+ 308 406 313 408 309 310 311 409 795 407 940 410 568 314 312 796 411 785 793 315
+ 316 792 317 318 941 413 302 787 791 319 799 414 320 412 650 415 35 801 797 651
+ 805 569 786 802 656 800
+ ICV_79 $T=0 0 0 0 $X=-25000 $Y=484000
X92 p_shift_out<1> VDDPST VDD VSS 39 322 917 25 324 333 323 280 335 332 918 327 328 325 326 331
+ 919 337 359 928 416 417 329 330 418 942 338 334 920 354 342 374 339 340 925 355
+ 341 371 336 898 346 923 922 357 817 343 900 345 364 924 837 419 347 348 349 27
+ 904 250 370 33 38 943 899 350 823 840 351 352 366 252 926 819 344 927 356 907
+ 169 830 360 921 353 388 383 363 362 365 930 361 367 376 929 368 369 378 373 358
+ 372 804 380 385 931 377 386 381 932 382 387 389 933 391 390 392 379 269 384 809
+ 934 393 394 395 790 397 935 401 398 938 937 936 396 399 409 408 403 402 415 939
+ 404 400 833 816 405 407 406 863 788 818 410 853 843 940 821 414 856 855 859 841
+ 824 847 860 842 839 941 850 851 807 825 811 852 827 814 411 822 857 413 37 861
+ 826 412 34 858 832 834 820 35 831 838 854 813 815 649 862 812 828 627 844 650
+ 36 849 848 808 864 835 845 829 810 648 846 806 664 836
+ ICV_78 $T=0 0 0 0 $X=-25000 $Y=597670
X93 p_shift_out<5> p_shift_out<6> VDDPST VSS VDD 25 39 942 943 ICV_73 $T=0 0 0 0 $X=-25000 $Y=743000
X94 VDDPST VDD VSS 27 25 39 p_shift_out<4> ICV_27 $T=0 210000 0 270 $X=0 $Y=129400
X95 VDDPST VDD VSS 25 129 39 p_shift_out<3> ICV_25 $T=0 290000 0 270 $X=0 $Y=209400
X96 VDDPST VSS ICV_23 $T=0 370000 0 270 $X=0 $Y=289400
X97 VDDPST VDD VSS ICV_18 $T=0 530000 0 270 $X=0 $Y=449400
X98 VDDPST VDD VSS 33 25 39 p_shift_out<2> ICV_11 $T=0 610000 0 270 $X=0 $Y=529400
X99 VDDPST VDD VSS 25 416 39 p_shift_out<0> ICV_9 $T=0 770000 0 270 $X=0 $Y=689400
X100 28 VSS VDD 717 128 421 728 420 118 112 722 726 439 723 725 714 724 713 423 435
+ 727 718 443 716 422 719 436 432 425 715 720 440 123 424 430 712 427 429 428 441
+ 426 721 437 944 431 433 434 438 945 442 444 445 446 947 466 946 451 448 447 450
+ 456 449 452 453 454 455 457 458 459 462 460 468 461 463 467 464 465 39 948 950
+ 470 469 473 490 486 471 479 487 484 952 472 478 476 482 480 477 949 951 481 475
+ 483 485 493 865 488 489 491 492
+ ICV_70 $T=0 0 0 0 $X=448710 $Y=154765
X101 30 VSS VDD 749 742 747 730 421 225 737 714 735 748 733 734 118 222 29 731 745
+ 126 432 420 494 750 495 739 740 741 422 510 216 729 214 425 123 423 736 498 499
+ 743 224 427 497 496 732 738 433 429 426 428 501 500 502 503 944 221 515 430 431
+ 505 434 112 946 953 508 962 506 507 509 552 961 436 444 964 438 511 437 435 951
+ 512 945 963 514 439 744 519 523 531 517 516 718 424 440 441 443 450 518 520 525
+ 954 597 457 446 521 453 524 522 447 445 526 448 449 466 452 947 451 530 513 533
+ 532 529 456 955 535 454 455 462 616 458 956 534 949 459 528 460 536 537 463 538
+ 461 746 504 539 541 464 950 465 540 958 467 468 959 470 527 542 544 551 543 471
+ 490 479 473 960 487 549 952 469 486 545 546 957 484 481 474 488 555 477 478 547
+ 548 553 557 475 476 550 554 480 866 558 556 482 965 485 483 559 560 491 492 561
+ 489
+ ICV_67 $T=0 0 0 0 $X=448710 $Y=241000
X102 VDD VSS VDDPST 775 217 755 763 777 780 31 758 753 756 771 318 779 496 759 764 774
+ 319 770 760 751 754 35 752 222 772 296 575 762 742 563 782 309 498 761 565 765
+ 32 564 494 221 776 783 953 781 567 768 568 757 773 569 566 570 769 571 497 778
+ 580 576 766 572 767 573 574 788 500 280 225 582 499 577 579 578 594 589 581 509
+ 501 584 503 970 592 966 505 271 502 504 585 586 525 587 26 544 604 588 518 506
+ 960 590 591 583 507 427 547 508 596 545 593 617 512 602 595 510 968 513 597 515
+ 530 519 517 520 598 954 269 599 521 948 609 524 514 608 516 600 601 523 603 534
+ 956 529 969 522 527 536 605 528 532 559 606 531 614 610 533 955 611 613 612 535
+ 957 607 615 538 620 616 540 511 618 959 958 537 539 619 703 624 622 972 542 541
+ 639 623 546 472 625 967 632 973 543 553 628 549 629 707 626 621 478 706 550 630
+ 634 558 627 631 633 555 635 636 950 551 962 638 554 637 804 557 548 971 645 951
+ 640 556 965 641 560 643 642 644 561
+ ICV_63 $T=0 0 0 0 $X=448710 $Y=358600
X103 VDD VSS 787 413 794 390 403 784 793 415 795 562 786 388 646 647 649 565 564 797
+ 35 650 563 572 566 788 803 789 357 798 571 648 404 785 585 321 796 659 570 800
+ 652 576 792 805 790 687 654 374 567 354 799 658 627 653 575 791 655 269 574 967
+ 694 577 579 525 581 662 801 580 802 804 573 660 582 583 584 586 663 966 664 637
+ 588 665 587 750 592 578 668 669 666 589 974 667 590 975 591 670 672 593 677 671
+ 680 676 657 594 595 674 596 656 597 547 661 599 978 685 673 969 675 601 598 976
+ 602 679 604 540 605 968 600 681 977 607 979 693 609 697 615 684 606 683 611 608
+ 603 682 983 686 688 613 612 614 678 980 981 526 539 696 617 622 689 690 619 985
+ 691 620 626 625 984 695 610 616 707 635 630 628 629 703 511 699 986 698 623 692
+ 631 632 633 634 973 636 987 945 706 961 700 702 704 951 701 552 963 962 638 705
+ 964 982 639 640 559 641 642 40 643 708 645 644
+ ICV_56 $T=0 0 0 0 $X=448710 $Y=484000
X104 p_shift_in<1> VDDPST VDD VSS 37 36 852 35 817 823 830 842 847 375 813 857 849 855 850 808
+ 835 843 809 861 399 836 841 834 837 854 862 851 839 788 821 826 810 846 820 647
+ 653 860 838 859 649 825 815 652 650 651 863 812 831 806 34 832 646 840 858 864
+ 818 845 819 848 811 828 853 654 824 709 655 816 827 814 636 822 657 656 844 660
+ 658 807 621 661 662 663 974 664 659 856 833 665 975 690 666 627 668 669 829 984
+ 670 667 671 618 643 676 674 677 678 673 680 686 977 976 681 675 978 970 682 979
+ 982 710 981 683 685 971 684 980 687 688 679 672 624 222 689 699 707 691 692 693
+ 695 694 983 696 623 697 945 985 972 628 698 986 703 632 804 706 987 961 700 701
+ 946 951 705 963 962 702 704 552 964 41 708 39 25
+ ICV_53 $T=0 0 0 0 $X=448710 $Y=597670
X105 VDD p_shift_in<7> p_shift_in<6> p_shift_in<5> VDDPST VSS 442 39 25 474 493 ICV_72 $T=0 0 0 0 $X=449000 $Y=-25000
X106 VDD p_shift_out<7> ack_p rstn_p VDDPST VSS 38 25 39 572 710 ICV_34 $T=0 0 0 0 $X=449000 $Y=743000
X107 VDDPST VDD VSS 39 25 865 p_shift_in<4> ICV_26 $T=900240 130000 0 90 $X=780240 $Y=129400
X108 VDDPST VDD VSS 39 25 866 p_shift_in<3> ICV_24 $T=900240 210000 0 90 $X=780240 $Y=209400
X109 VDDPST VSS ICV_22 $T=900240 290000 0 90 $X=780240 $Y=289400
X110 VDDPST VDD VSS ICV_17 $T=900240 450000 0 90 $X=780240 $Y=449400
X111 VDDPST VDD VSS 40 39 25 p_shift_in<2> ICV_10 $T=900240 530000 0 90 $X=780240 $Y=529400
X112 VDDPST VDD VSS 39 41 25 p_shift_in<0> ICV_8 $T=900240 690000 0 90 $X=780240 $Y=689400
.ENDS
***************************************
