* SPICE NETLIST
***************************************

.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT mimcap_1p0_sin TOP BOT
.ENDS
***************************************
.SUBCKT mimcap_1p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin TOP BOT
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT na20_g5a_cfp_mac D G S B
.ENDS
***************************************
.SUBCKT na20_g5a_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT na29_g5a_cfp_mac D G S B
.ENDS
***************************************
.SUBCKT na29_g5a_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT na6_g5a_nbl_v2_mac D G S B SUB
.ENDS
***************************************
.SUBCKT nch_hv5_5vnw_ac D G S B
.ENDS
***************************************
.SUBCKT nda29_g3a_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT nda45_g3b_nbl_cfp_mac D G BS SUB
.ENDS
***************************************
.SUBCKT ndio_sbd_mac PLUS MINUS
.ENDS
***************************************
.SUBCKT nld12_g5a_cfp_mac D G BS
.ENDS
***************************************
.SUBCKT nld12_g5a_iso_cfp_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld16_g5a_cfp_mac D G BS
.ENDS
***************************************
.SUBCKT nld16_g5a_iso_cfp_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld20_g5a_cfp_mac D G BS
.ENDS
***************************************
.SUBCKT nld20_g5a_iso_cfp_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld24_g5a_cfp_mac D G BS
.ENDS
***************************************
.SUBCKT nld24_g5a_iso_cfp_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld24_g5a_iso_switch_cfp_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld24_g5a_switch_cfp_mac D G BS
.ENDS
***************************************
.SUBCKT nld36_g5b_nbl_cfp_mac D G BS SUB
.ENDS
***************************************
.SUBCKT nld45_g5b_nbl_cfp_mac D G BS SUB
.ENDS
***************************************
.SUBCKT nld5_g5a_iso_switch_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld6_g5a_de_iso_v2_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld6_g5a_de_mac D G BS
.ENDS
***************************************
.SUBCKT nld6_g5a_sa_iso_v2_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld6_g5a_sa_mac D G BS
.ENDS
***************************************
.SUBCKT nld9_g5a_iso_mac D G BS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nld9_g5a_mac D G BS
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_5 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_5_mis PLUS MINUS
.ENDS
***************************************
.SUBCKT npddshnnbl10_ga_bgr8_7t C1 C8 B1 B8 E1 E8 SUB
.ENDS
***************************************
.SUBCKT npddshnnbl10_ga_poly_4t C B E SUB
.ENDS
***************************************
.SUBCKT npddshnnbl2_ga_poly_4t C B E SUB
.ENDS
***************************************
.SUBCKT npddshnnbl5_ga_poly_4t C B E SUB
.ENDS
***************************************
.SUBCKT npwshnnbl10_ga_bgr8_7t C1 C8 B1 B8 E1 E8 SUB
.ENDS
***************************************
.SUBCKT npwshnnbl10_ga_poly_4t C B E SUB
.ENDS
***************************************
.SUBCKT npwshnnbl2_ga_poly_4t C B E SUB
.ENDS
***************************************
.SUBCKT npwshnnbl5_ga_poly_4t C B E SUB
.ENDS
***************************************
.SUBCKT pa12_g5a_nbl_slit_v2_mac D G BS SUB
.ENDS
***************************************
.SUBCKT pa12_g5a_nbl_v2_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa16_g5a_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa16_g5a_nbl_slit_cfp_mac D G BS SUB
.ENDS
***************************************
.SUBCKT pa20_g5a_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa20_g5a_nbl_slit_cfp_mac D G BS SUB
.ENDS
***************************************
.SUBCKT pa29_g5a_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa36_g5b_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa45_g5b_nbl_cfp_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa6_g5a_de_nbl_v2_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa6_g5a_sa_nbl_v2_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa9_g5a_nbl_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pa9_g5a_nbl_slit_mac D G BS SUB
.ENDS
***************************************
.SUBCKT pbhvnwshnnbl_esd_dio_shp_gb_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pbshnnbl_dio_shp_ga_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pch5_as_switch_mac D G BS SUB
.ENDS
***************************************
.SUBCKT pddshnnbl_dio_shp_ga_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_12_pdd_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_12_v4_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_16_v3_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_20_pdd_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_20_v3_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_24_v3_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_29_v3_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_6_v3_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_ga_9_v3_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_gb_36_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pdio_esd_gb_45_cit_v3_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT phvnwpsub10_gb_poly C B E
.ENDS
***************************************
.SUBCKT phvnwpsub2_gb_poly C B E
.ENDS
***************************************
.SUBCKT phvnwpsub5_gb_poly C B E
.ENDS
***************************************
.SUBCKT pnddpsub10_ga_poly C B E
.ENDS
***************************************
.SUBCKT pnddpsub2_ga_poly C B E
.ENDS
***************************************
.SUBCKT pnddpsub5_ga_poly C B E
.ENDS
***************************************
.SUBCKT pnddshp5_nbl_ga_4t C B E SUB
.ENDS
***************************************
.SUBCKT rnod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodrpo_pure5v PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodrpo_pure5v_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1rpo_pure5v PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpo1rpo_pure5v_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwod_pure5v PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_pure5v_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwsti_pure5v PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_pure5v_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodrpo_pure5v PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodrpo_pure5v_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1rpo_pure5v PLUS MINUS
.ENDS
***************************************
.SUBCKT rppo1rpo_pure5v_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1rpo_serp PLUS MINUS
.ENDS
***************************************
.SUBCKT rppo1rpo_serp_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppolyhri1k PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyhri1k_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyhri3d3k PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyhri3d3k_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyhri3d3k_serp PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyhri3d3k_serp_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_dio_ga_12_v2_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT sbd_dio_ga_16_v2_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT sbd_dio_ga_24_v2_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT shpnblshn_dio_shp_gb_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT shpshnnbl_esd_dio_shp_ga_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT zd_dio_ga_nbl_v2_4t PLUS MINUS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT TAPCELLBWP7T
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ANTENNABWP7T VSS I
** N=3 EP=2 IP=0 FDC=1
D0 VSS I DN AREA=2.037e-13 PJ=1.81e-06 $X=140 $Y=520 $D=32
.ENDS
***************************************
.SUBCKT ICV_1 1 3 4
** N=4 EP=3 IP=6 FDC=2
X0 1 3 ANTENNABWP7T $T=0 0 0 0 $X=-290 $Y=-235
X1 1 4 ANTENNABWP7T $T=1120 0 0 0 $X=830 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_2 1 3 4
** N=4 EP=3 IP=6 FDC=2
X0 1 3 ANTENNABWP7T $T=-1120 0 0 0 $X=-1410 $Y=-235
X1 1 4 ANTENNABWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT FILL1BWP7T
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CKBD1BWP7T I VSS VDD Z
** N=5 EP=4 IP=0 FDC=4
M0 VSS I 5 VSS N L=1.8e-07 W=4.55e-07 $X=620 $Y=425 $D=0
M1 Z 5 VSS VSS N L=1.8e-07 W=5.2e-07 $X=1440 $Y=360 $D=0
M2 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M3 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1440 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INVD0BWP7T I VSS VDD ZN
** N=4 EP=4 IP=0 FDC=2
M0 ZN I VSS VSS N L=1.8e-07 W=5e-07 $X=840 $Y=560 $D=0
M1 ZN I VDD VDD P L=1.8e-07 W=6.85e-07 $X=840 $Y=2575 $D=16
.ENDS
***************************************
.SUBCKT BUFFD1P5BWP7T I Z VSS VDD
** N=5 EP=4 IP=0 FDC=6
M0 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 VSS 5 Z VSS N L=1.8e-07 W=4.65e-07 $X=2060 $Y=880 $D=0
M3 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M4 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M5 VDD 5 Z VDD P L=1.8e-07 W=6.85e-07 $X=2060 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INVD3BWP7T I VSS VDD ZN
** N=4 EP=4 IP=0 FDC=6
M0 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=885 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=1605 $Y=345 $D=0
M2 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=2535 $Y=345 $D=0
M3 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=885 $Y=2205 $D=16
M4 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1605 $Y=2205 $D=16
M5 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=2535 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT MAOI22D0BWP7T B1 B2 VDD VSS A1 ZN A2
** N=11 EP=7 IP=0 FDC=10
M0 8 B1 VSS VSS N L=1.8e-07 W=5e-07 $X=460 $Y=845 $D=0
M1 VSS B2 8 VSS N L=1.8e-07 W=5e-07 $X=1180 $Y=845 $D=0
M2 ZN 8 VSS VSS N L=1.8e-07 W=5e-07 $X=1980 $Y=845 $D=0
M3 9 A1 ZN VSS N L=1.8e-07 W=5e-07 $X=2700 $Y=845 $D=0
M4 VSS A2 9 VSS N L=1.8e-07 W=5e-07 $X=3280 $Y=845 $D=0
M5 10 B1 8 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2625 $D=16
M6 VDD B2 10 VDD P L=1.8e-07 W=6.85e-07 $X=1050 $Y=2625 $D=16
M7 11 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1850 $Y=2625 $D=16
M8 ZN A1 11 VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2300 $D=16
M9 11 A2 ZN VDD P L=1.8e-07 W=6.85e-07 $X=3280 $Y=2300 $D=16
.ENDS
***************************************
.SUBCKT FILL2BWP7T
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MAOI22D2BWP7T A1 A2 B1 B2 ZN VSS VDD
** N=12 EP=7 IP=0 FDC=14
M0 11 A1 8 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS A2 11 VSS N L=1.8e-07 W=1e-06 $X=1060 $Y=345 $D=0
M2 9 8 VSS VSS N L=1.8e-07 W=1e-06 $X=1780 $Y=345 $D=0
M3 10 B1 9 VSS N L=1.8e-07 W=1e-06 $X=2500 $Y=345 $D=0
M4 9 B2 10 VSS N L=1.8e-07 W=1e-06 $X=3220 $Y=345 $D=0
M5 ZN 10 VSS VSS N L=1.8e-07 W=1e-06 $X=4640 $Y=345 $D=0
M6 VSS 10 ZN VSS N L=1.8e-07 W=1e-06 $X=5360 $Y=345 $D=0
M7 8 A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M8 VDD A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M9 10 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M10 12 B1 10 VDD P L=1.8e-07 W=1.37e-06 $X=2785 $Y=2205 $D=16
M11 VDD B2 12 VDD P L=1.8e-07 W=1.37e-06 $X=3380 $Y=2205 $D=16
M12 ZN 10 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4640 $Y=2205 $D=16
M13 VDD 10 ZN VDD P L=1.8e-07 W=1.37e-06 $X=5360 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IAO22D2BWP7T A2 A1 ZN B1 VSS B2 VDD
** N=12 EP=7 IP=0 FDC=14
M0 8 10 9 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS A2 8 VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 8 A1 VSS VSS N L=1.8e-07 W=1e-06 $X=2140 $Y=345 $D=0
M3 ZN 9 VSS VSS N L=1.8e-07 W=1e-06 $X=3490 $Y=345 $D=0
M4 VSS 9 ZN VSS N L=1.8e-07 W=1e-06 $X=4210 $Y=345 $D=0
M5 11 B1 VSS VSS N L=1.8e-07 W=5e-07 $X=4930 $Y=345 $D=0
M6 10 B2 11 VSS N L=1.8e-07 W=5e-07 $X=5360 $Y=345 $D=0
M7 9 10 VDD VDD P L=1.8e-07 W=1.37e-06 $X=685 $Y=2205 $D=16
M8 12 A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=1405 $Y=2205 $D=16
M9 VDD A1 12 VDD P L=1.8e-07 W=1.37e-06 $X=1965 $Y=2205 $D=16
M10 ZN 9 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2795 $Y=2205 $D=16
M11 VDD 9 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3840 $Y=2205 $D=16
M12 10 B1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=4640 $Y=2820 $D=16
M13 VDD B2 10 VDD P L=1.8e-07 W=6.85e-07 $X=5360 $Y=2820 $D=16
.ENDS
***************************************
.SUBCKT BUFFD1BWP7T I VSS VDD Z
** N=5 EP=4 IP=0 FDC=4
M0 VSS I 5 VSS N L=1.8e-07 W=5e-07 $X=625 $Y=845 $D=0
M1 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=1425 $Y=345 $D=0
M2 VDD I 5 VDD P L=1.8e-07 W=6.85e-07 $X=625 $Y=2205 $D=16
M3 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1425 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT DCAP4BWP7T VSS VDD
** N=4 EP=2 IP=0 FDC=4
M0 VSS 4 VSS VSS N L=2.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 3 4 VSS VSS N L=1.8e-07 W=1e-06 $X=1440 $Y=345 $D=0
M2 VDD 3 VDD VDD P L=2.8e-07 W=1.17e-06 $X=620 $Y=2405 $D=16
M3 4 3 VDD VDD P L=1.8e-07 W=1.17e-06 $X=1440 $Y=2405 $D=16
.ENDS
***************************************
.SUBCKT ICV_3 1 2
** N=2 EP=2 IP=4 FDC=4
X1 1 2 DCAP4BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT DCAP8BWP7T VSS VDD
** N=4 EP=2 IP=0 FDC=6
M0 VSS 4 VSS VSS N L=9.9e-07 W=9.45e-07 $X=620 $Y=345 $D=0
M1 VSS 4 VSS VSS N L=9.9e-07 W=9.45e-07 $X=2150 $Y=345 $D=0
M2 3 4 VSS VSS N L=1.8e-07 W=9.45e-07 $X=3680 $Y=345 $D=0
M3 VDD 3 VDD VDD P L=9.9e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M4 VDD 3 VDD VDD P L=9.9e-07 W=1.235e-06 $X=2150 $Y=2340 $D=16
M5 4 3 VDD VDD P L=1.8e-07 W=1.235e-06 $X=3680 $Y=2340 $D=16
.ENDS
***************************************
.SUBCKT DCAPBWP7T VDD VSS
** N=4 EP=2 IP=0 FDC=2
M0 3 4 VSS VSS N L=1.8e-07 W=1e-06 $X=800 $Y=345 $D=0
M1 4 3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=680 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AO222D0BWP7T B2 A1 A2 B1 C1 C2 VSS VDD Z
** N=15 EP=9 IP=0 FDC=14
M0 12 A1 11 VSS N L=1.8e-07 W=5e-07 $X=1085 $Y=455 $D=0
M1 VSS A2 12 VSS N L=1.8e-07 W=5e-07 $X=1555 $Y=455 $D=0
M2 13 B2 VSS VSS N L=1.8e-07 W=5e-07 $X=2355 $Y=455 $D=0
M3 11 B1 13 VSS N L=1.8e-07 W=5e-07 $X=2825 $Y=455 $D=0
M4 14 C1 11 VSS N L=1.8e-07 W=5e-07 $X=3615 $Y=455 $D=0
M5 VSS C2 14 VSS N L=1.8e-07 W=5e-07 $X=4250 $Y=455 $D=0
M6 Z 11 VSS VSS N L=1.8e-07 W=5e-07 $X=5360 $Y=455 $D=0
M7 15 B2 10 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2760 $D=16
M8 11 A1 15 VDD P L=1.8e-07 W=6.85e-07 $X=1240 $Y=2500 $D=16
M9 15 A2 11 VDD P L=1.8e-07 W=6.85e-07 $X=1960 $Y=2500 $D=16
M10 10 B1 15 VDD P L=1.8e-07 W=6.85e-07 $X=2580 $Y=2500 $D=16
M11 VDD C1 10 VDD P L=1.8e-07 W=6.85e-07 $X=3300 $Y=2500 $D=16
M12 10 C2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=4100 $Y=2500 $D=16
M13 Z 11 VDD VDD P L=1.8e-07 W=6.85e-07 $X=5360 $Y=2300 $D=16
.ENDS
***************************************
.SUBCKT OAI221D1BWP7T C VSS B2 B1 A2 VDD ZN A1
** N=12 EP=8 IP=0 FDC=10
M0 9 C VSS VSS N L=1.8e-07 W=1e-06 $X=625 $Y=345 $D=0
M1 10 B2 9 VSS N L=1.8e-07 W=1e-06 $X=1345 $Y=345 $D=0
M2 9 B1 10 VSS N L=1.8e-07 W=1e-06 $X=2065 $Y=345 $D=0
M3 ZN A2 10 VSS N L=1.8e-07 W=1e-06 $X=3520 $Y=345 $D=0
M4 10 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=4240 $Y=345 $D=0
M5 ZN C VDD VDD P L=1.8e-07 W=1.37e-06 $X=625 $Y=2205 $D=16
M6 11 B2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1345 $Y=2205 $D=16
M7 VDD B1 11 VDD P L=1.8e-07 W=1.37e-06 $X=1825 $Y=2205 $D=16
M8 12 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3520 $Y=2205 $D=16
M9 ZN A1 12 VDD P L=1.8e-07 W=1.37e-06 $X=4240 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AO222D1BWP7T A2 A1 B1 B2 C1 C2 VSS VDD Z
** N=15 EP=9 IP=0 FDC=14
M0 13 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 12 A1 13 VSS N L=1.8e-07 W=1e-06 $X=1345 $Y=345 $D=0
M2 14 B1 12 VSS N L=1.8e-07 W=1e-06 $X=2065 $Y=345 $D=0
M3 VSS B2 14 VSS N L=1.8e-07 W=1e-06 $X=2580 $Y=345 $D=0
M4 15 C1 12 VSS N L=1.8e-07 W=1e-06 $X=4300 $Y=345 $D=0
M5 VSS C2 15 VSS N L=1.8e-07 W=1e-06 $X=5020 $Y=345 $D=0
M6 Z 12 VSS VSS N L=1.8e-07 W=1e-06 $X=5920 $Y=345 $D=0
M7 12 A2 10 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M8 10 A1 12 VDD P L=1.8e-07 W=1.37e-06 $X=1345 $Y=2205 $D=16
M9 11 B1 10 VDD P L=1.8e-07 W=1.37e-06 $X=2065 $Y=2205 $D=16
M10 10 B2 11 VDD P L=1.8e-07 W=1.37e-06 $X=2840 $Y=2205 $D=16
M11 11 C1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4300 $Y=2205 $D=16
M12 VDD C2 11 VDD P L=1.8e-07 W=1.37e-06 $X=5020 $Y=2205 $D=16
M13 Z 12 VDD VDD P L=1.8e-07 W=1.37e-06 $X=5920 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_4 1 2
** N=2 EP=2 IP=4 FDC=6
X0 1 2 DCAP4BWP7T $T=0 0 0 0 $X=-290 $Y=-235
X1 2 1 DCAPBWP7T $T=2240 0 0 0 $X=1950 $Y=-235
.ENDS
***************************************
.SUBCKT DFCNQD1BWP7T CP D CDN VDD VSS Q
** N=19 EP=6 IP=0 FDC=28
M0 VSS CP 7 VSS N L=1.8e-07 W=5e-07 $X=640 $Y=840 $D=0
M1 8 7 VSS VSS N L=1.8e-07 W=5e-07 $X=1240 $Y=840 $D=0
M2 15 7 VSS VSS N L=1.8e-07 W=9.4e-07 $X=2660 $Y=405 $D=0
M3 10 D 15 VSS N L=1.8e-07 W=9.4e-07 $X=3160 $Y=405 $D=0
M4 16 8 10 VSS N L=1.8e-07 W=4.2e-07 $X=4005 $Y=895 $D=0
M5 17 CDN 16 VSS N L=1.8e-07 W=4.2e-07 $X=4435 $Y=895 $D=0
M6 VSS 11 17 VSS N L=1.8e-07 W=4.2e-07 $X=4865 $Y=895 $D=0
M7 11 10 VSS VSS N L=1.8e-07 W=5.4e-07 $X=5715 $Y=775 $D=0
M8 13 8 11 VSS N L=1.8e-07 W=9.1e-07 $X=6435 $Y=405 $D=0
M9 12 7 13 VSS N L=1.8e-07 W=4.2e-07 $X=7255 $Y=895 $D=0
M10 VSS 14 12 VSS N L=1.8e-07 W=4.2e-07 $X=8915 $Y=895 $D=0
M11 18 CDN VSS VSS N L=1.8e-07 W=9.7e-07 $X=9610 $Y=345 $D=0
M12 14 13 18 VSS N L=1.8e-07 W=9.7e-07 $X=10055 $Y=345 $D=0
M13 Q 14 VSS VSS N L=1.8e-07 W=1e-06 $X=11520 $Y=345 $D=0
M14 VDD CP 7 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2345 $D=16
M15 8 7 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1240 $Y=2345 $D=16
M16 19 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2525 $Y=2205 $D=16
M17 10 D 19 VDD P L=1.8e-07 W=1.37e-06 $X=2955 $Y=2205 $D=16
M18 9 7 10 VDD P L=1.8e-07 W=4.2e-07 $X=3795 $Y=2365 $D=16
M19 VDD CDN 9 VDD P L=1.8e-07 W=4.2e-07 $X=4515 $Y=2365 $D=16
M20 9 11 VDD VDD P L=1.8e-07 W=4.2e-07 $X=5115 $Y=2365 $D=16
M21 11 10 VDD VDD P L=1.8e-07 W=6.2e-07 $X=6375 $Y=2175 $D=16
M22 13 7 11 VDD P L=1.8e-07 W=6.2e-07 $X=7255 $Y=2175 $D=16
M23 12 8 13 VDD P L=1.8e-07 W=4.2e-07 $X=8080 $Y=2175 $D=16
M24 VDD 14 12 VDD P L=1.8e-07 W=4.2e-07 $X=8915 $Y=2175 $D=16
M25 14 CDN VDD VDD P L=1.8e-07 W=4.2e-07 $X=9850 $Y=3095 $D=16
M26 VDD 13 14 VDD P L=1.8e-07 W=1.37e-06 $X=10680 $Y=2205 $D=16
M27 Q 14 VDD VDD P L=1.8e-07 W=1.37e-06 $X=11520 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_5
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT FILL16BWP7T
** N=19 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILL8BWP7T
** N=11 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILL4BWP7T
** N=7 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_8 1 2
** N=2 EP=2 IP=4 FDC=4
X1 1 2 ICV_3 $T=1120 0 0 0 $X=830 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_9 1 2
** N=2 EP=2 IP=4 FDC=6
X1 1 2 DCAP8BWP7T $T=1120 0 0 0 $X=830 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_10 1 2
** N=2 EP=2 IP=4 FDC=4
X1 1 2 DCAP4BWP7T $T=1120 0 0 0 $X=830 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_11
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13 1 2
** N=2 EP=2 IP=4 FDC=4
X1 1 2 DCAP4BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT MAOI22D1BWP7T B1 B2 VDD A1 ZN A2 VSS
** N=11 EP=7 IP=0 FDC=10
M0 8 B1 VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS B2 8 VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 ZN 8 VSS VSS N L=1.8e-07 W=1e-06 $X=2150 $Y=345 $D=0
M3 10 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=2955 $Y=345 $D=0
M4 VSS A2 10 VSS N L=1.8e-07 W=1e-06 $X=3680 $Y=345 $D=0
M5 11 B1 8 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M6 VDD B2 11 VDD P L=1.8e-07 W=1.37e-06 $X=1330 $Y=2205 $D=16
M7 9 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2150 $Y=2205 $D=16
M8 ZN A1 9 VDD P L=1.8e-07 W=1.37e-06 $X=2955 $Y=2205 $D=16
M9 9 A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3680 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IOA21D0BWP7T A1 A2 VSS ZN B VDD
** N=9 EP=6 IP=0 FDC=8
M0 8 A1 7 VSS N L=1.8e-07 W=4.2e-07 $X=625 $Y=440 $D=0
M1 VSS A2 8 VSS N L=1.8e-07 W=4.2e-07 $X=1205 $Y=440 $D=0
M2 9 7 VSS VSS N L=1.8e-07 W=5e-07 $X=1945 $Y=360 $D=0
M3 ZN B 9 VSS N L=1.8e-07 W=5e-07 $X=2560 $Y=360 $D=0
M4 7 A1 VDD VDD P L=1.8e-07 W=4.2e-07 $X=465 $Y=2500 $D=16
M5 VDD A2 7 VDD P L=1.8e-07 W=4.2e-07 $X=1185 $Y=2500 $D=16
M6 ZN 7 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1840 $Y=2500 $D=16
M7 VDD B ZN VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2500 $D=16
.ENDS
***************************************
.SUBCKT INVD1BWP7T I VSS VDD ZN
** N=4 EP=4 IP=0 FDC=2
M0 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=840 $Y=345 $D=0
M1 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=840 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_14 1 2
** N=2 EP=2 IP=4 FDC=6
X1 1 2 DCAP8BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=34
X0 1 2 DCAP8BWP7T $T=0 0 1 180 $X=-4770 $Y=-235
X1 3 4 5 2 1 6 DFCNQD1BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT BUFFD10BWP7T I Z VSS VDD
** N=5 EP=4 IP=0 FDC=28
M0 5 I VSS VSS N L=1.8e-07 W=4.65e-07 $X=460 $Y=880 $D=0
M1 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=1180 $Y=345 $D=0
M2 5 I VSS VSS N L=1.8e-07 W=1e-06 $X=1900 $Y=345 $D=0
M3 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=2620 $Y=345 $D=0
M4 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=3340 $Y=345 $D=0
M5 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=4060 $Y=345 $D=0
M6 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=4780 $Y=345 $D=0
M7 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=5500 $Y=345 $D=0
M8 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=6220 $Y=345 $D=0
M9 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=6940 $Y=345 $D=0
M10 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=7660 $Y=345 $D=0
M11 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=8380 $Y=345 $D=0
M12 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=9120 $Y=345 $D=0
M13 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=9840 $Y=345 $D=0
M14 5 I VDD VDD P L=1.8e-07 W=8.35e-07 $X=460 $Y=2205 $D=16
M15 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=1180 $Y=2205 $D=16
M16 5 I VDD VDD P L=1.8e-07 W=1.37e-06 $X=1900 $Y=2205 $D=16
M17 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=2620 $Y=2205 $D=16
M18 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3340 $Y=2205 $D=16
M19 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=4060 $Y=2205 $D=16
M20 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4780 $Y=2205 $D=16
M21 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=5500 $Y=2205 $D=16
M22 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=6220 $Y=2205 $D=16
M23 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=6940 $Y=2205 $D=16
M24 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=7660 $Y=2205 $D=16
M25 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=8380 $Y=2205 $D=16
M26 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=9120 $Y=2205 $D=16
M27 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=9840 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT BUFFD2BWP7T I Z VSS VDD
** N=5 EP=4 IP=0 FDC=6
M0 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=680 $Y=345 $D=0
M1 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=1590 $Y=345 $D=0
M2 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=2430 $Y=345 $D=0
M3 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=680 $Y=2205 $D=16
M4 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1590 $Y=2205 $D=16
M5 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=2430 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT DFCNQD2BWP7T CP D CDN Q VSS VDD
** N=19 EP=6 IP=0 FDC=30
M0 VSS CP 7 VSS N L=1.8e-07 W=5e-07 $X=640 $Y=840 $D=0
M1 8 7 VSS VSS N L=1.8e-07 W=5e-07 $X=1240 $Y=840 $D=0
M2 15 7 VSS VSS N L=1.8e-07 W=9.4e-07 $X=2660 $Y=405 $D=0
M3 10 D 15 VSS N L=1.8e-07 W=9.4e-07 $X=3160 $Y=405 $D=0
M4 16 8 10 VSS N L=1.8e-07 W=4.2e-07 $X=4005 $Y=895 $D=0
M5 17 CDN 16 VSS N L=1.8e-07 W=4.2e-07 $X=4435 $Y=895 $D=0
M6 VSS 11 17 VSS N L=1.8e-07 W=4.2e-07 $X=4865 $Y=895 $D=0
M7 11 10 VSS VSS N L=1.8e-07 W=5.4e-07 $X=5715 $Y=775 $D=0
M8 13 8 11 VSS N L=1.8e-07 W=9.1e-07 $X=6435 $Y=405 $D=0
M9 12 7 13 VSS N L=1.8e-07 W=4.2e-07 $X=7200 $Y=895 $D=0
M10 VSS 14 12 VSS N L=1.8e-07 W=4.2e-07 $X=8910 $Y=895 $D=0
M11 18 CDN VSS VSS N L=1.8e-07 W=9.7e-07 $X=9510 $Y=345 $D=0
M12 14 13 18 VSS N L=1.8e-07 W=9.7e-07 $X=9940 $Y=345 $D=0
M13 Q 14 VSS VSS N L=1.8e-07 W=1e-06 $X=11360 $Y=345 $D=0
M14 VSS 14 Q VSS N L=1.8e-07 W=1e-06 $X=12080 $Y=345 $D=0
M15 VDD CP 7 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2345 $D=16
M16 8 7 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1240 $Y=2345 $D=16
M17 19 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2525 $Y=2205 $D=16
M18 10 D 19 VDD P L=1.8e-07 W=1.37e-06 $X=2955 $Y=2205 $D=16
M19 9 7 10 VDD P L=1.8e-07 W=4.2e-07 $X=3795 $Y=2365 $D=16
M20 VDD CDN 9 VDD P L=1.8e-07 W=4.2e-07 $X=4515 $Y=2365 $D=16
M21 9 11 VDD VDD P L=1.8e-07 W=4.2e-07 $X=5115 $Y=2365 $D=16
M22 11 10 VDD VDD P L=1.8e-07 W=6.2e-07 $X=6375 $Y=2175 $D=16
M23 13 7 11 VDD P L=1.8e-07 W=6.2e-07 $X=7300 $Y=2175 $D=16
M24 12 8 13 VDD P L=1.8e-07 W=4.2e-07 $X=8115 $Y=2175 $D=16
M25 VDD 14 12 VDD P L=1.8e-07 W=4.2e-07 $X=8895 $Y=2175 $D=16
M26 14 CDN VDD VDD P L=1.8e-07 W=4.2e-07 $X=9850 $Y=3095 $D=16
M27 VDD 13 14 VDD P L=1.8e-07 W=1.37e-06 $X=10630 $Y=2205 $D=16
M28 Q 14 VDD VDD P L=1.8e-07 W=1.37e-06 $X=11360 $Y=2205 $D=16
M29 VDD 14 Q VDD P L=1.8e-07 W=1.37e-06 $X=12080 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT DCAP16BWP7T VSS VDD
** N=4 EP=2 IP=0 FDC=12
M0 VSS 4 VSS VSS N L=9.65e-07 W=9.4e-07 $X=620 $Y=405 $D=0
M1 VSS 4 VSS VSS N L=9.65e-07 W=9.4e-07 $X=2125 $Y=405 $D=0
M2 VSS 4 VSS VSS N L=9.65e-07 W=9.4e-07 $X=3630 $Y=405 $D=0
M3 VSS 4 VSS VSS N L=9.65e-07 W=9.4e-07 $X=5135 $Y=405 $D=0
M4 VSS 4 VSS VSS N L=9.65e-07 W=9.4e-07 $X=6640 $Y=405 $D=0
M5 3 4 VSS VSS N L=1.8e-07 W=9.4e-07 $X=8160 $Y=405 $D=0
M6 VDD 3 VDD VDD P L=9.65e-07 W=1.31e-06 $X=620 $Y=2205 $D=16
M7 VDD 3 VDD VDD P L=9.65e-07 W=1.31e-06 $X=2125 $Y=2205 $D=16
M8 VDD 3 VDD VDD P L=9.65e-07 W=1.31e-06 $X=3630 $Y=2205 $D=16
M9 VDD 3 VDD VDD P L=9.65e-07 W=1.31e-06 $X=5135 $Y=2205 $D=16
M10 VDD 3 VDD VDD P L=9.65e-07 W=1.095e-06 $X=6640 $Y=2420 $D=16
M11 4 3 VDD VDD P L=1.8e-07 W=1.095e-06 $X=8160 $Y=2420 $D=16
.ENDS
***************************************
.SUBCKT CKND1BWP7T I VSS VDD ZN
** N=4 EP=4 IP=0 FDC=2
M0 ZN I VSS VSS N L=1.8e-07 W=5.25e-07 $X=830 $Y=440 $D=0
M1 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=830 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INVD4BWP7T I ZN VSS VDD
** N=4 EP=4 IP=0 FDC=8
M0 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=765 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=1485 $Y=345 $D=0
M2 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=2275 $Y=345 $D=0
M3 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=2995 $Y=345 $D=0
M4 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=765 $Y=2205 $D=16
M5 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1485 $Y=2205 $D=16
M6 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=2275 $Y=2205 $D=16
M7 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=2995 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT BUFFD3BWP7T I VSS VDD Z
** N=5 EP=4 IP=0 FDC=8
M0 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=680 $Y=345 $D=0
M1 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=1570 $Y=345 $D=0
M2 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=2400 $Y=345 $D=0
M3 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=3120 $Y=345 $D=0
M4 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=680 $Y=2205 $D=16
M5 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1570 $Y=2205 $D=16
M6 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=2400 $Y=2205 $D=16
M7 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3120 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT BUFFD12BWP7T I Z VSS VDD
** N=5 EP=4 IP=0 FDC=32
M0 5 I VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 5 I VSS VSS N L=1.8e-07 W=1e-06 $X=2060 $Y=345 $D=0
M3 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=2780 $Y=345 $D=0
M4 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=3500 $Y=345 $D=0
M5 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=4220 $Y=345 $D=0
M6 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=4940 $Y=345 $D=0
M7 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=5660 $Y=345 $D=0
M8 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=6400 $Y=345 $D=0
M9 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=7120 $Y=345 $D=0
M10 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=7850 $Y=345 $D=0
M11 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=8570 $Y=345 $D=0
M12 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=9300 $Y=345 $D=0
M13 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=10020 $Y=345 $D=0
M14 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=10740 $Y=345 $D=0
M15 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=11500 $Y=345 $D=0
M16 5 I VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M17 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M18 5 I VDD VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M19 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M20 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3500 $Y=2205 $D=16
M21 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=4220 $Y=2205 $D=16
M22 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4940 $Y=2205 $D=16
M23 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=5660 $Y=2205 $D=16
M24 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=6400 $Y=2205 $D=16
M25 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=7120 $Y=2205 $D=16
M26 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=7850 $Y=2205 $D=16
M27 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=8570 $Y=2205 $D=16
M28 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=9300 $Y=2205 $D=16
M29 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=10020 $Y=2205 $D=16
M30 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=10740 $Y=2205 $D=16
M31 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=11500 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKXOR2D4BWP7T A1 A2 Z VSS VDD
** N=9 EP=5 IP=0 FDC=27
M0 7 8 VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=570 $D=0
M1 VSS 8 7 VSS N L=1.8e-07 W=5e-07 $X=1340 $Y=570 $D=0
M2 6 A1 VSS VSS N L=1.8e-07 W=5.25e-07 $X=2210 $Y=545 $D=0
M3 7 A1 9 VSS N L=1.8e-07 W=4.2e-07 $X=3780 $Y=830 $D=0
M4 9 A1 7 VSS N L=1.8e-07 W=4.2e-07 $X=4500 $Y=830 $D=0
M5 8 6 9 VSS N L=1.8e-07 W=4.2e-07 $X=5220 $Y=830 $D=0
M6 9 6 8 VSS N L=1.8e-07 W=4.2e-07 $X=5940 $Y=830 $D=0
M7 8 A2 VSS VSS N L=1.8e-07 W=7.5e-07 $X=7640 $Y=555 $D=0
M8 VSS A2 8 VSS N L=1.8e-07 W=7.5e-07 $X=8420 $Y=555 $D=0
M9 Z 9 VSS VSS N L=1.8e-07 W=6e-07 $X=9360 $Y=555 $D=0
M10 VSS 9 Z VSS N L=1.8e-07 W=6e-07 $X=10080 $Y=555 $D=0
M11 Z 9 VSS VSS N L=1.8e-07 W=6e-07 $X=10800 $Y=555 $D=0
M12 VSS 9 Z VSS N L=1.8e-07 W=6e-07 $X=11520 $Y=555 $D=0
M13 7 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M14 VDD 8 7 VDD P L=1.8e-07 W=1.645e-06 $X=1340 $Y=1930 $D=16
M15 6 A1 VDD VDD P L=1.8e-07 W=1.31e-06 $X=2180 $Y=2110 $D=16
M16 7 6 9 VDD P L=1.8e-07 W=1.035e-06 $X=3620 $Y=2110 $D=16
M17 9 6 7 VDD P L=1.8e-07 W=1.035e-06 $X=4340 $Y=2110 $D=16
M18 8 A1 9 VDD P L=1.8e-07 W=1.13e-06 $X=5060 $Y=2370 $D=16
M19 9 A1 8 VDD P L=1.8e-07 W=1.13e-06 $X=5780 $Y=2370 $D=16
M20 VDD A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=7200 $Y=2205 $D=16
M21 8 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=7920 $Y=2205 $D=16
M22 VDD A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=8640 $Y=2205 $D=16
M23 Z 9 VDD VDD P L=1.8e-07 W=1.37e-06 $X=9360 $Y=2205 $D=16
M24 VDD 9 Z VDD P L=1.8e-07 W=1.37e-06 $X=10080 $Y=2205 $D=16
M25 Z 9 VDD VDD P L=1.8e-07 W=1.37e-06 $X=10800 $Y=2205 $D=16
M26 VDD 9 Z VDD P L=1.8e-07 W=1.37e-06 $X=11520 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AOI22D1BWP7T B1 B2 VDD A2 VSS A1 ZN
** N=10 EP=7 IP=0 FDC=8
M0 9 B1 ZN VSS N L=1.8e-07 W=1e-06 $X=640 $Y=345 $D=0
M1 VSS B2 9 VSS N L=1.8e-07 W=1e-06 $X=1440 $Y=345 $D=0
M2 10 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=2420 $Y=345 $D=0
M3 ZN A1 10 VSS N L=1.8e-07 W=1e-06 $X=3120 $Y=345 $D=0
M4 VDD B1 8 VDD P L=1.8e-07 W=1.37e-06 $X=640 $Y=2205 $D=16
M5 8 B2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1440 $Y=2205 $D=16
M6 ZN A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=2180 $Y=2205 $D=16
M7 8 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3120 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OAI21D1BWP7T A1 A2 VDD B ZN VSS
** N=8 EP=6 IP=0 FDC=6
M0 ZN A1 7 VSS N L=1.8e-07 W=1e-06 $X=760 $Y=345 $D=0
M1 7 A2 ZN VSS N L=1.8e-07 W=1e-06 $X=1480 $Y=345 $D=0
M2 VSS B 7 VSS N L=1.8e-07 W=1e-06 $X=2200 $Y=345 $D=0
M3 8 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=760 $Y=2205 $D=16
M4 VDD A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=1480 $Y=2205 $D=16
M5 ZN B VDD VDD P L=1.8e-07 W=1.37e-06 $X=2200 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKND12BWP7T I VDD ZN VSS
** N=4 EP=4 IP=0 FDC=22
M0 ZN I VSS VSS N L=1.8e-07 W=6.3e-07 $X=1340 $Y=410 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=6.3e-07 $X=2060 $Y=410 $D=0
M2 ZN I VSS VSS N L=1.8e-07 W=6.3e-07 $X=2780 $Y=410 $D=0
M3 VSS I ZN VSS N L=1.8e-07 W=6.3e-07 $X=3500 $Y=410 $D=0
M4 ZN I VSS VSS N L=1.8e-07 W=6.3e-07 $X=4220 $Y=410 $D=0
M5 VSS I ZN VSS N L=1.8e-07 W=6.3e-07 $X=4940 $Y=410 $D=0
M6 ZN I VSS VSS N L=1.8e-07 W=6.3e-07 $X=5660 $Y=410 $D=0
M7 VSS I ZN VSS N L=1.8e-07 W=6.3e-07 $X=6380 $Y=410 $D=0
M8 ZN I VSS VSS N L=1.8e-07 W=6.3e-07 $X=7100 $Y=410 $D=0
M9 VSS I ZN VSS N L=1.8e-07 W=6.3e-07 $X=7820 $Y=410 $D=0
M10 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M11 VDD I ZN VDD P L=1.8e-07 W=1.525e-06 $X=1340 $Y=2050 $D=16
M12 ZN I VDD VDD P L=1.8e-07 W=1.525e-06 $X=2060 $Y=2050 $D=16
M13 VDD I ZN VDD P L=1.8e-07 W=1.525e-06 $X=2780 $Y=2050 $D=16
M14 ZN I VDD VDD P L=1.8e-07 W=1.525e-06 $X=3500 $Y=2050 $D=16
M15 VDD I ZN VDD P L=1.8e-07 W=1.525e-06 $X=4220 $Y=2050 $D=16
M16 ZN I VDD VDD P L=1.8e-07 W=1.525e-06 $X=4940 $Y=2050 $D=16
M17 VDD I ZN VDD P L=1.8e-07 W=1.525e-06 $X=5660 $Y=2050 $D=16
M18 ZN I VDD VDD P L=1.8e-07 W=1.525e-06 $X=6380 $Y=2050 $D=16
M19 VDD I ZN VDD P L=1.8e-07 W=1.525e-06 $X=7100 $Y=2050 $D=16
M20 ZN I VDD VDD P L=1.8e-07 W=1.345e-06 $X=7820 $Y=2230 $D=16
D21 VSS I DN AREA=2.037e-13 PJ=1.81e-06 $X=140 $Y=645 $D=32
.ENDS
***************************************
.SUBCKT BUFFD8BWP7T I Z VSS VDD
** N=5 EP=4 IP=0 FDC=22
M0 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 5 I VSS VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=2060 $Y=345 $D=0
M3 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=2780 $Y=345 $D=0
M4 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=3500 $Y=345 $D=0
M5 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=4220 $Y=345 $D=0
M6 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=4940 $Y=345 $D=0
M7 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=5660 $Y=345 $D=0
M8 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=6380 $Y=345 $D=0
M9 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=7100 $Y=345 $D=0
M10 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=7820 $Y=345 $D=0
M11 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M12 5 I VDD VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M13 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M14 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M15 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=3500 $Y=2205 $D=16
M16 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4220 $Y=2205 $D=16
M17 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=4940 $Y=2205 $D=16
M18 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=5660 $Y=2205 $D=16
M19 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=6380 $Y=2205 $D=16
M20 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=7100 $Y=2205 $D=16
M21 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=7820 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR2D4BWP7T A2 VDD A1 ZN VSS
** N=6 EP=5 IP=0 FDC=16
M0 ZN A2 VSS VSS N L=1.8e-07 W=1e-06 $X=660 $Y=345 $D=0
M1 VSS A2 ZN VSS N L=1.8e-07 W=1e-06 $X=1380 $Y=345 $D=0
M2 ZN A2 VSS VSS N L=1.8e-07 W=1e-06 $X=2100 $Y=345 $D=0
M3 VSS A2 ZN VSS N L=1.8e-07 W=1e-06 $X=2820 $Y=345 $D=0
M4 ZN A1 VSS VSS N L=1.8e-07 W=1e-06 $X=3540 $Y=345 $D=0
M5 VSS A1 ZN VSS N L=1.8e-07 W=1e-06 $X=4260 $Y=345 $D=0
M6 ZN A1 VSS VSS N L=1.8e-07 W=1e-06 $X=4980 $Y=345 $D=0
M7 VSS A1 ZN VSS N L=1.8e-07 W=1e-06 $X=5700 $Y=345 $D=0
M8 VDD A2 6 VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M9 6 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1380 $Y=2205 $D=16
M10 VDD A2 6 VDD P L=1.8e-07 W=1.37e-06 $X=2100 $Y=2205 $D=16
M11 6 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2820 $Y=2205 $D=16
M12 ZN A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=3540 $Y=2205 $D=16
M13 6 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4260 $Y=2205 $D=16
M14 ZN A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=4980 $Y=2205 $D=16
M15 6 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=5700 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AO21D0BWP7T A2 A1 B VSS VDD Z
** N=9 EP=6 IP=0 FDC=8
M0 8 A2 VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=460 $D=0
M1 7 A1 8 VSS N L=1.8e-07 W=5e-07 $X=1120 $Y=460 $D=0
M2 VSS B 7 VSS N L=1.8e-07 W=5e-07 $X=1840 $Y=460 $D=0
M3 Z 7 VSS VSS N L=1.8e-07 W=5e-07 $X=2560 $Y=460 $D=0
M4 7 A2 9 VDD P L=1.8e-07 W=6.85e-07 $X=490 $Y=2555 $D=16
M5 9 A1 7 VDD P L=1.8e-07 W=6.85e-07 $X=1210 $Y=2555 $D=16
M6 VDD B 9 VDD P L=1.8e-07 W=6.85e-07 $X=1840 $Y=2555 $D=16
M7 Z 7 VDD VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2555 $D=16
.ENDS
***************************************
.SUBCKT BUFFD6BWP7T I Z VSS VDD
** N=5 EP=4 IP=0 FDC=16
M0 5 I VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=2080 $Y=345 $D=0
M3 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=2800 $Y=345 $D=0
M4 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=3520 $Y=345 $D=0
M5 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=4240 $Y=345 $D=0
M6 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=4960 $Y=345 $D=0
M7 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=5680 $Y=345 $D=0
M8 5 I VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M9 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M10 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2080 $Y=2205 $D=16
M11 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=2800 $Y=2205 $D=16
M12 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3520 $Y=2205 $D=16
M13 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=4240 $Y=2205 $D=16
M14 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4960 $Y=2205 $D=16
M15 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=5680 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INVD2BWP7T I ZN VDD VSS
** N=4 EP=4 IP=0 FDC=4
M0 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=670 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=1390 $Y=345 $D=0
M2 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=670 $Y=2205 $D=16
M3 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1390 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKXOR2D1BWP7T A1 A2 VSS VDD Z
** N=10 EP=5 IP=0 FDC=12
M0 VSS A1 6 VSS N L=1.8e-07 W=9.4e-07 $X=620 $Y=405 $D=0
M1 9 7 VSS VSS N L=1.8e-07 W=4.2e-07 $X=1380 $Y=830 $D=0
M2 8 A1 9 VSS N L=1.8e-07 W=4.2e-07 $X=1980 $Y=440 $D=0
M3 7 6 8 VSS N L=1.8e-07 W=4.2e-07 $X=2740 $Y=830 $D=0
M4 VSS A2 7 VSS N L=1.8e-07 W=4.2e-07 $X=3520 $Y=440 $D=0
M5 Z 8 VSS VSS N L=1.8e-07 W=8e-07 $X=4240 $Y=440 $D=0
M6 VDD A1 6 VDD P L=1.8e-07 W=6e-07 $X=620 $Y=2205 $D=16
M7 10 7 VDD VDD P L=1.8e-07 W=9.4e-07 $X=1420 $Y=2205 $D=16
M8 8 6 10 VDD P L=1.8e-07 W=9.4e-07 $X=1960 $Y=2205 $D=16
M9 7 A1 8 VDD P L=1.8e-07 W=1.185e-06 $X=2690 $Y=2205 $D=16
M10 VDD A2 7 VDD P L=1.8e-07 W=1e-06 $X=3480 $Y=2205 $D=16
M11 Z 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4240 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKXOR2D2BWP7T A1 A2 Z VSS VDD
** N=10 EP=5 IP=0 FDC=14
M0 VSS A1 6 VSS N L=1.8e-07 W=9.4e-07 $X=620 $Y=405 $D=0
M1 9 7 VSS VSS N L=1.8e-07 W=4.2e-07 $X=1380 $Y=775 $D=0
M2 8 A1 9 VSS N L=1.8e-07 W=6e-07 $X=1980 $Y=405 $D=0
M3 7 6 8 VSS N L=1.8e-07 W=8e-07 $X=2780 $Y=450 $D=0
M4 VSS A2 7 VSS N L=1.8e-07 W=6e-07 $X=3795 $Y=450 $D=0
M5 Z 8 VSS VSS N L=1.8e-07 W=1e-06 $X=4600 $Y=345 $D=0
M6 VSS 8 Z VSS N L=1.8e-07 W=1e-06 $X=5320 $Y=345 $D=0
M7 VDD A1 6 VDD P L=1.8e-07 W=6e-07 $X=620 $Y=2205 $D=16
M8 10 7 VDD VDD P L=1.8e-07 W=1.2e-06 $X=1420 $Y=2375 $D=16
M9 8 6 10 VDD P L=1.8e-07 W=1.2e-06 $X=1960 $Y=2375 $D=16
M10 7 A1 8 VDD P L=1.8e-07 W=1.185e-06 $X=2780 $Y=2375 $D=16
M11 VDD A2 7 VDD P L=1.8e-07 W=1.2e-06 $X=3800 $Y=2375 $D=16
M12 Z 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4600 $Y=2205 $D=16
M13 VDD 8 Z VDD P L=1.8e-07 W=1.37e-06 $X=5320 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT DCAP32BWP7T VDD VSS
** N=4 EP=2 IP=0 FDC=24
M0 VSS 3 4 VSS N L=1.8e-07 W=9.4e-07 $X=620 $Y=405 $D=0
M1 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=1340 $Y=405 $D=0
M2 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=2915 $Y=405 $D=0
M3 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=4490 $Y=405 $D=0
M4 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=6065 $Y=405 $D=0
M5 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=7640 $Y=405 $D=0
M6 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=9215 $Y=405 $D=0
M7 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=10790 $Y=405 $D=0
M8 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=12365 $Y=405 $D=0
M9 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=13940 $Y=405 $D=0
M10 VSS 3 VSS VSS N L=1.035e-06 W=9.4e-07 $X=15515 $Y=405 $D=0
M11 4 3 VSS VSS N L=1.8e-07 W=9.4e-07 $X=17120 $Y=405 $D=0
M12 VDD 4 3 VDD P L=1.8e-07 W=1.095e-06 $X=620 $Y=2420 $D=16
M13 VDD 4 VDD VDD P L=1.035e-06 W=1.095e-06 $X=1340 $Y=2420 $D=16
M14 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=2915 $Y=2205 $D=16
M15 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=4490 $Y=2205 $D=16
M16 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=6065 $Y=2205 $D=16
M17 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=7640 $Y=2205 $D=16
M18 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=9215 $Y=2205 $D=16
M19 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=10790 $Y=2205 $D=16
M20 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=12365 $Y=2205 $D=16
M21 VDD 4 VDD VDD P L=1.035e-06 W=1.31e-06 $X=13940 $Y=2205 $D=16
M22 VDD 4 VDD VDD P L=1.035e-06 W=1.095e-06 $X=15515 $Y=2420 $D=16
M23 3 4 VDD VDD P L=1.8e-07 W=1.095e-06 $X=17120 $Y=2420 $D=16
.ENDS
***************************************
.SUBCKT XNR4D1BWP7T A4 A3 ZN A2 A1 VSS VDD
** N=21 EP=7 IP=0 FDC=30
M0 VSS A4 8 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=500 $D=0
M1 16 9 VSS VSS N L=1.8e-07 W=5e-07 $X=1445 $Y=845 $D=0
M2 10 A4 16 VSS N L=1.8e-07 W=5e-07 $X=1925 $Y=845 $D=0
M3 9 8 10 VSS N L=1.8e-07 W=5e-07 $X=2645 $Y=845 $D=0
M4 VSS A3 9 VSS N L=1.8e-07 W=1e-06 $X=3425 $Y=345 $D=0
M5 VSS 10 11 VSS N L=1.8e-07 W=5e-07 $X=4980 $Y=775 $D=0
M6 17 13 VSS VSS N L=1.8e-07 W=5e-07 $X=5700 $Y=775 $D=0
M7 12 10 17 VSS N L=1.8e-07 W=5e-07 $X=6180 $Y=775 $D=0
M8 13 11 12 VSS N L=1.8e-07 W=5e-07 $X=6900 $Y=775 $D=0
M9 VSS 12 ZN VSS N L=1.8e-07 W=1e-06 $X=8320 $Y=345 $D=0
M10 14 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=9120 $Y=345 $D=0
M11 13 15 14 VSS N L=1.8e-07 W=5e-07 $X=9885 $Y=775 $D=0
M12 18 A1 13 VSS N L=1.8e-07 W=5e-07 $X=10605 $Y=775 $D=0
M13 VSS 14 18 VSS N L=1.8e-07 W=5e-07 $X=11320 $Y=775 $D=0
M14 15 A1 VSS VSS N L=1.8e-07 W=5e-07 $X=12080 $Y=595 $D=0
M15 VDD A4 8 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2710 $D=16
M16 19 9 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1380 $Y=2460 $D=16
M17 10 8 19 VDD P L=1.8e-07 W=6.85e-07 $X=1925 $Y=2460 $D=16
M18 9 A4 10 VDD P L=1.8e-07 W=6.85e-07 $X=2645 $Y=2460 $D=16
M19 VDD A3 9 VDD P L=1.8e-07 W=1.37e-06 $X=3425 $Y=2205 $D=16
M20 VDD 10 11 VDD P L=1.8e-07 W=6.85e-07 $X=4980 $Y=2370 $D=16
M21 20 13 VDD VDD P L=1.8e-07 W=6.85e-07 $X=5700 $Y=2370 $D=16
M22 12 11 20 VDD P L=1.8e-07 W=6.85e-07 $X=6180 $Y=2370 $D=16
M23 13 10 12 VDD P L=1.8e-07 W=6.85e-07 $X=6900 $Y=2370 $D=16
M24 VDD 12 ZN VDD P L=1.8e-07 W=1.31e-06 $X=8320 $Y=2205 $D=16
M25 14 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=9120 $Y=2205 $D=16
M26 13 A1 14 VDD P L=1.8e-07 W=6.85e-07 $X=9885 $Y=2385 $D=16
M27 21 15 13 VDD P L=1.8e-07 W=6.85e-07 $X=10605 $Y=2385 $D=16
M28 VDD 14 21 VDD P L=1.8e-07 W=6.85e-07 $X=11290 $Y=2385 $D=16
M29 15 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=12080 $Y=2720 $D=16
.ENDS
***************************************
.SUBCKT BUFFD5BWP7T I VSS VDD Z
** N=5 EP=4 IP=0 FDC=14
M0 5 I VSS VSS N L=1.8e-07 W=1e-06 $X=640 $Y=345 $D=0
M1 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=1360 $Y=345 $D=0
M2 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=2140 $Y=345 $D=0
M3 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=2860 $Y=345 $D=0
M4 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=3640 $Y=345 $D=0
M5 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=4360 $Y=345 $D=0
M6 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=5140 $Y=345 $D=0
M7 5 I VDD VDD P L=1.8e-07 W=1.37e-06 $X=640 $Y=2205 $D=16
M8 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=1360 $Y=2205 $D=16
M9 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2140 $Y=2205 $D=16
M10 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=2860 $Y=2205 $D=16
M11 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3640 $Y=2205 $D=16
M12 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=4360 $Y=2205 $D=16
M13 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=5140 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OAI21D0BWP7T A2 ZN A1 B VSS VDD
** N=8 EP=6 IP=0 FDC=6
M0 ZN A2 7 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=845 $D=0
M1 7 A1 ZN VSS N L=1.8e-07 W=5e-07 $X=1340 $Y=845 $D=0
M2 VSS B 7 VSS N L=1.8e-07 W=4.65e-07 $X=2060 $Y=880 $D=0
M3 8 A2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2770 $D=16
M4 ZN A1 8 VDD P L=1.8e-07 W=6.85e-07 $X=1250 $Y=2770 $D=16
M5 VDD B ZN VDD P L=1.8e-07 W=6.85e-07 $X=1975 $Y=2770 $D=16
.ENDS
***************************************
.SUBCKT XNR4D0BWP7T A4 A3 ZN A2 A1 VSS VDD
** N=21 EP=7 IP=0 FDC=30
M0 VSS A4 8 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=500 $D=0
M1 16 9 VSS VSS N L=1.8e-07 W=5e-07 $X=1445 $Y=835 $D=0
M2 10 A4 16 VSS N L=1.8e-07 W=5e-07 $X=1925 $Y=835 $D=0
M3 9 8 10 VSS N L=1.8e-07 W=5e-07 $X=2645 $Y=835 $D=0
M4 VSS A3 9 VSS N L=1.8e-07 W=5e-07 $X=3425 $Y=835 $D=0
M5 VSS 10 11 VSS N L=1.8e-07 W=5e-07 $X=4980 $Y=775 $D=0
M6 17 13 VSS VSS N L=1.8e-07 W=5e-07 $X=5700 $Y=775 $D=0
M7 12 10 17 VSS N L=1.8e-07 W=5e-07 $X=6180 $Y=775 $D=0
M8 13 11 12 VSS N L=1.8e-07 W=5e-07 $X=6900 $Y=775 $D=0
M9 VSS 12 ZN VSS N L=1.8e-07 W=5e-07 $X=8320 $Y=630 $D=0
M10 14 A2 VSS VSS N L=1.8e-07 W=5e-07 $X=9120 $Y=630 $D=0
M11 13 15 14 VSS N L=1.8e-07 W=5e-07 $X=9885 $Y=775 $D=0
M12 18 A1 13 VSS N L=1.8e-07 W=5e-07 $X=10605 $Y=775 $D=0
M13 VSS 14 18 VSS N L=1.8e-07 W=5e-07 $X=11320 $Y=775 $D=0
M14 15 A1 VSS VSS N L=1.8e-07 W=5e-07 $X=12080 $Y=595 $D=0
M15 VDD A4 8 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2710 $D=16
M16 19 9 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1380 $Y=2460 $D=16
M17 10 8 19 VDD P L=1.8e-07 W=6.85e-07 $X=1925 $Y=2460 $D=16
M18 9 A4 10 VDD P L=1.8e-07 W=6.85e-07 $X=2645 $Y=2460 $D=16
M19 VDD A3 9 VDD P L=1.8e-07 W=6.85e-07 $X=3425 $Y=2205 $D=16
M20 VDD 10 11 VDD P L=1.8e-07 W=6.85e-07 $X=4980 $Y=2370 $D=16
M21 20 13 VDD VDD P L=1.8e-07 W=6.85e-07 $X=5700 $Y=2370 $D=16
M22 12 11 20 VDD P L=1.8e-07 W=6.85e-07 $X=6180 $Y=2370 $D=16
M23 13 10 12 VDD P L=1.8e-07 W=6.85e-07 $X=6900 $Y=2370 $D=16
M24 VDD 12 ZN VDD P L=1.8e-07 W=6.85e-07 $X=8320 $Y=2205 $D=16
M25 14 A2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=9120 $Y=2205 $D=16
M26 13 A1 14 VDD P L=1.8e-07 W=6.85e-07 $X=9885 $Y=2385 $D=16
M27 21 15 13 VDD P L=1.8e-07 W=6.85e-07 $X=10605 $Y=2385 $D=16
M28 VDD 14 21 VDD P L=1.8e-07 W=6.85e-07 $X=11290 $Y=2385 $D=16
M29 15 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=12080 $Y=2720 $D=16
.ENDS
***************************************
.SUBCKT XNR4D2BWP7T A4 A3 ZN A2 A1 VSS VDD
** N=21 EP=7 IP=0 FDC=32
M0 VSS A4 8 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=500 $D=0
M1 16 9 VSS VSS N L=1.8e-07 W=5e-07 $X=1445 $Y=845 $D=0
M2 10 A4 16 VSS N L=1.8e-07 W=5e-07 $X=1925 $Y=845 $D=0
M3 9 8 10 VSS N L=1.8e-07 W=5e-07 $X=2645 $Y=845 $D=0
M4 VSS A3 9 VSS N L=1.8e-07 W=1e-06 $X=3425 $Y=345 $D=0
M5 VSS 10 11 VSS N L=1.8e-07 W=5e-07 $X=4980 $Y=775 $D=0
M6 17 13 VSS VSS N L=1.8e-07 W=5e-07 $X=5700 $Y=775 $D=0
M7 12 10 17 VSS N L=1.8e-07 W=5e-07 $X=6180 $Y=775 $D=0
M8 13 11 12 VSS N L=1.8e-07 W=5e-07 $X=6900 $Y=775 $D=0
M9 ZN 12 VSS VSS N L=1.8e-07 W=1e-06 $X=8320 $Y=345 $D=0
M10 VSS 12 ZN VSS N L=1.8e-07 W=1e-06 $X=9040 $Y=345 $D=0
M11 14 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=9800 $Y=345 $D=0
M12 13 15 14 VSS N L=1.8e-07 W=5e-07 $X=10580 $Y=775 $D=0
M13 18 A1 13 VSS N L=1.8e-07 W=5e-07 $X=11300 $Y=775 $D=0
M14 VSS 14 18 VSS N L=1.8e-07 W=5e-07 $X=11880 $Y=775 $D=0
M15 15 A1 VSS VSS N L=1.8e-07 W=5e-07 $X=12640 $Y=595 $D=0
M16 VDD A4 8 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2710 $D=16
M17 19 9 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1380 $Y=2460 $D=16
M18 10 8 19 VDD P L=1.8e-07 W=6.85e-07 $X=1925 $Y=2460 $D=16
M19 9 A4 10 VDD P L=1.8e-07 W=6.85e-07 $X=2645 $Y=2460 $D=16
M20 VDD A3 9 VDD P L=1.8e-07 W=1.37e-06 $X=3425 $Y=2205 $D=16
M21 VDD 10 11 VDD P L=1.8e-07 W=6.85e-07 $X=4980 $Y=2370 $D=16
M22 20 13 VDD VDD P L=1.8e-07 W=6.85e-07 $X=5700 $Y=2370 $D=16
M23 12 11 20 VDD P L=1.8e-07 W=6.85e-07 $X=6180 $Y=2370 $D=16
M24 13 10 12 VDD P L=1.8e-07 W=6.85e-07 $X=6900 $Y=2370 $D=16
M25 ZN 12 VDD VDD P L=1.8e-07 W=1.37e-06 $X=8320 $Y=2205 $D=16
M26 VDD 12 ZN VDD P L=1.8e-07 W=1.37e-06 $X=9040 $Y=2205 $D=16
M27 14 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=9800 $Y=2205 $D=16
M28 13 A1 14 VDD P L=1.8e-07 W=6.85e-07 $X=10580 $Y=2385 $D=16
M29 21 15 13 VDD P L=1.8e-07 W=6.85e-07 $X=11300 $Y=2385 $D=16
M30 VDD 14 21 VDD P L=1.8e-07 W=6.85e-07 $X=11880 $Y=2385 $D=16
M31 15 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=12640 $Y=2720 $D=16
.ENDS
***************************************
.SUBCKT MUX2ND1BWP7T I0 S I1 VSS VDD ZN
** N=13 EP=6 IP=0 FDC=14
M0 VSS S 7 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=345 $D=0
M1 10 I0 VSS VSS N L=1.8e-07 W=1e-06 $X=1375 $Y=345 $D=0
M2 8 7 10 VSS N L=1.8e-07 W=5e-07 $X=1980 $Y=345 $D=0
M3 11 S 8 VSS N L=1.8e-07 W=5e-07 $X=2700 $Y=345 $D=0
M4 VSS I1 11 VSS N L=1.8e-07 W=1e-06 $X=3310 $Y=345 $D=0
M5 9 8 VSS VSS N L=1.8e-07 W=5e-07 $X=4030 $Y=345 $D=0
M6 ZN 9 VSS VSS N L=1.8e-07 W=1e-06 $X=5360 $Y=345 $D=0
M7 VDD S 7 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2590 $D=16
M8 12 I0 VDD VDD P L=1.8e-07 W=9.4e-07 $X=1385 $Y=2205 $D=16
M9 8 S 12 VDD P L=1.8e-07 W=6.85e-07 $X=1990 $Y=2590 $D=16
M10 13 7 8 VDD P L=1.8e-07 W=6.85e-07 $X=2710 $Y=2590 $D=16
M11 VDD I1 13 VDD P L=1.8e-07 W=1.37e-06 $X=3310 $Y=2205 $D=16
M12 9 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=4030 $Y=2580 $D=16
M13 ZN 9 VDD VDD P L=1.8e-07 W=1.37e-06 $X=5360 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT XNR3D2BWP7T A2 A1 A3 ZN VSS VDD
** N=16 EP=6 IP=0 FDC=24
M0 VSS A2 7 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=500 $D=0
M1 13 8 VSS VSS N L=1.8e-07 W=5e-07 $X=1380 $Y=845 $D=0
M2 9 7 13 VSS N L=1.8e-07 W=5e-07 $X=1840 $Y=845 $D=0
M3 8 A2 9 VSS N L=1.8e-07 W=5e-07 $X=2600 $Y=715 $D=0
M4 VSS A1 8 VSS N L=1.8e-07 W=1e-06 $X=3320 $Y=345 $D=0
M5 VSS 9 10 VSS N L=1.8e-07 W=6.4e-07 $X=4770 $Y=705 $D=0
M6 14 11 VSS VSS N L=1.8e-07 W=5.7e-07 $X=5530 $Y=775 $D=0
M7 12 10 14 VSS N L=1.8e-07 W=5.7e-07 $X=6200 $Y=775 $D=0
M8 11 9 12 VSS N L=1.8e-07 W=5e-07 $X=6920 $Y=845 $D=0
M9 VSS A3 11 VSS N L=1.8e-07 W=1e-06 $X=7665 $Y=345 $D=0
M10 ZN 12 VSS VSS N L=1.8e-07 W=1e-06 $X=8560 $Y=345 $D=0
M11 VSS 12 ZN VSS N L=1.8e-07 W=1e-06 $X=9280 $Y=345 $D=0
M12 VDD A2 7 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2205 $D=16
M13 15 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1380 $Y=2205 $D=16
M14 9 A2 15 VDD P L=1.8e-07 W=6.85e-07 $X=1980 $Y=2335 $D=16
M15 8 7 9 VDD P L=1.8e-07 W=6.85e-07 $X=2700 $Y=2205 $D=16
M16 VDD A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=3420 $Y=2205 $D=16
M17 VDD 9 10 VDD P L=1.8e-07 W=8.25e-07 $X=4770 $Y=2205 $D=16
M18 16 11 VDD VDD P L=1.8e-07 W=9.35e-07 $X=5530 $Y=2205 $D=16
M19 12 9 16 VDD P L=1.8e-07 W=8e-07 $X=6190 $Y=2410 $D=16
M20 11 10 12 VDD P L=1.8e-07 W=8.65e-07 $X=6910 $Y=2345 $D=16
M21 VDD A3 11 VDD P L=1.8e-07 W=1.37e-06 $X=7665 $Y=2205 $D=16
M22 ZN 12 VDD VDD P L=1.8e-07 W=1.37e-06 $X=8560 $Y=2205 $D=16
M23 VDD 12 ZN VDD P L=1.8e-07 W=1.37e-06 $X=9280 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT XNR2D1BWP7T A1 A2 VSS VDD ZN
** N=10 EP=5 IP=0 FDC=12
M0 VSS A1 6 VSS N L=1.8e-07 W=5e-07 $X=625 $Y=460 $D=0
M1 9 7 VSS VSS N L=1.8e-07 W=5e-07 $X=1425 $Y=845 $D=0
M2 8 6 9 VSS N L=1.8e-07 W=5e-07 $X=1855 $Y=845 $D=0
M3 7 A1 8 VSS N L=1.8e-07 W=5e-07 $X=2725 $Y=440 $D=0
M4 VSS A2 7 VSS N L=1.8e-07 W=1e-06 $X=3485 $Y=345 $D=0
M5 ZN 8 VSS VSS N L=1.8e-07 W=1e-06 $X=4235 $Y=345 $D=0
M6 VDD A1 6 VDD P L=1.8e-07 W=6.85e-07 $X=625 $Y=2530 $D=16
M7 10 7 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1425 $Y=2445 $D=16
M8 8 A1 10 VDD P L=1.8e-07 W=6.85e-07 $X=1935 $Y=2445 $D=16
M9 7 6 8 VDD P L=1.8e-07 W=6.85e-07 $X=2685 $Y=2445 $D=16
M10 VDD A2 7 VDD P L=1.8e-07 W=1.37e-06 $X=3465 $Y=2205 $D=16
M11 ZN 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4235 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKND2BWP7T I ZN VDD VSS
** N=4 EP=4 IP=0 FDC=4
M0 ZN I VSS VSS N L=1.8e-07 W=5.25e-07 $X=670 $Y=440 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=5.25e-07 $X=1390 $Y=440 $D=0
M2 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=670 $Y=2205 $D=16
M3 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1390 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKND0BWP7T I VSS VDD ZN
** N=4 EP=4 IP=0 FDC=2
M0 ZN I VSS VSS N L=1.8e-07 W=4.2e-07 $X=830 $Y=505 $D=0
M1 ZN I VDD VDD P L=1.8e-07 W=1.13e-06 $X=830 $Y=2445 $D=16
.ENDS
***************************************
.SUBCKT CKXOR2D0BWP7T A1 A2 VSS VDD Z
** N=10 EP=5 IP=0 FDC=12
M0 VSS A1 6 VSS N L=1.8e-07 W=9.4e-07 $X=620 $Y=405 $D=0
M1 9 7 VSS VSS N L=1.8e-07 W=4.2e-07 $X=1380 $Y=790 $D=0
M2 8 A1 9 VSS N L=1.8e-07 W=4.2e-07 $X=1980 $Y=440 $D=0
M3 7 6 8 VSS N L=1.8e-07 W=4.2e-07 $X=2740 $Y=830 $D=0
M4 VSS A2 7 VSS N L=1.8e-07 W=4.2e-07 $X=3520 $Y=440 $D=0
M5 Z 8 VSS VSS N L=1.8e-07 W=4.2e-07 $X=4240 $Y=440 $D=0
M6 VDD A1 6 VDD P L=1.8e-07 W=6e-07 $X=620 $Y=2205 $D=16
M7 10 7 VDD VDD P L=1.8e-07 W=9.4e-07 $X=1420 $Y=2205 $D=16
M8 8 6 10 VDD P L=1.8e-07 W=9.4e-07 $X=1960 $Y=2205 $D=16
M9 7 A1 8 VDD P L=1.8e-07 W=1.185e-06 $X=2690 $Y=2205 $D=16
M10 VDD A2 7 VDD P L=1.8e-07 W=9.4e-07 $X=3520 $Y=2620 $D=16
M11 Z 8 VDD VDD P L=1.8e-07 W=8.8e-07 $X=4240 $Y=2680 $D=16
.ENDS
***************************************
.SUBCKT IAO22D1BWP7T A2 A1 ZN B1 B2 VDD VSS
** N=11 EP=7 IP=0 FDC=10
M0 8 A2 VSS VSS N L=1.8e-07 W=7.7e-07 $X=665 $Y=575 $D=0
M1 VSS A1 8 VSS N L=1.8e-07 W=7.7e-07 $X=1425 $Y=575 $D=0
M2 ZN 8 VSS VSS N L=1.8e-07 W=1e-06 $X=2600 $Y=345 $D=0
M3 10 B1 ZN VSS N L=1.8e-07 W=1e-06 $X=3500 $Y=345 $D=0
M4 VSS B2 10 VSS N L=1.8e-07 W=1e-06 $X=4240 $Y=345 $D=0
M5 11 A2 VDD VDD P L=1.8e-07 W=1.17e-06 $X=665 $Y=2400 $D=16
M6 8 A1 11 VDD P L=1.8e-07 W=1.17e-06 $X=1265 $Y=2400 $D=16
M7 9 8 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2800 $Y=2205 $D=16
M8 VDD B1 9 VDD P L=1.8e-07 W=1.37e-06 $X=3520 $Y=2205 $D=16
M9 9 B2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4240 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AOI22D2BWP7T B1 VDD B2 ZN A1 A2 VSS
** N=12 EP=7 IP=0 FDC=16
M0 9 B2 VSS VSS N L=1.8e-07 W=1e-06 $X=630 $Y=345 $D=0
M1 ZN B1 9 VSS N L=1.8e-07 W=1e-06 $X=1400 $Y=345 $D=0
M2 10 B1 ZN VSS N L=1.8e-07 W=1e-06 $X=2120 $Y=345 $D=0
M3 VSS B2 10 VSS N L=1.8e-07 W=1e-06 $X=2760 $Y=345 $D=0
M4 11 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=3720 $Y=345 $D=0
M5 ZN A1 11 VSS N L=1.8e-07 W=1e-06 $X=4380 $Y=345 $D=0
M6 12 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=5140 $Y=345 $D=0
M7 VSS A2 12 VSS N L=1.8e-07 W=1e-06 $X=5680 $Y=345 $D=0
M8 VDD B2 8 VDD P L=1.8e-07 W=1.37e-06 $X=630 $Y=2205 $D=16
M9 8 B1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1400 $Y=2205 $D=16
M10 VDD B1 8 VDD P L=1.8e-07 W=1.37e-06 $X=2120 $Y=2205 $D=16
M11 8 B2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2880 $Y=2205 $D=16
M12 ZN A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=3640 $Y=2205 $D=16
M13 8 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4380 $Y=2205 $D=16
M14 ZN A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=5140 $Y=2205 $D=16
M15 8 A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=5860 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT MUX2ND0BWP7T S I0 I1 ZN VSS VDD
** N=11 EP=6 IP=0 FDC=10
M0 VSS S 7 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=345 $D=0
M1 8 I0 VSS VSS N L=1.8e-07 W=1e-06 $X=1385 $Y=345 $D=0
M2 ZN 7 8 VSS N L=1.8e-07 W=5e-07 $X=2005 $Y=345 $D=0
M3 9 S ZN VSS N L=1.8e-07 W=5e-07 $X=2725 $Y=345 $D=0
M4 VSS I1 9 VSS N L=1.8e-07 W=1e-06 $X=3535 $Y=345 $D=0
M5 VDD S 7 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2700 $D=16
M6 10 I0 VDD VDD P L=1.8e-07 W=9.4e-07 $X=1385 $Y=2205 $D=16
M7 ZN S 10 VDD P L=1.8e-07 W=6.85e-07 $X=2005 $Y=2590 $D=16
M8 11 7 ZN VDD P L=1.8e-07 W=6.85e-07 $X=2805 $Y=2590 $D=16
M9 VDD I1 11 VDD P L=1.8e-07 W=1.37e-06 $X=3535 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AOI22D0BWP7T B2 ZN A1 B1 A2 VDD VSS
** N=10 EP=7 IP=0 FDC=8
M0 8 B2 VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=345 $D=0
M1 ZN B1 8 VSS N L=1.8e-07 W=5e-07 $X=1165 $Y=345 $D=0
M2 9 A1 ZN VSS N L=1.8e-07 W=5e-07 $X=1940 $Y=345 $D=0
M3 VSS A2 9 VSS N L=1.8e-07 W=5e-07 $X=2560 $Y=345 $D=0
M4 10 B2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2755 $D=16
M5 ZN A1 10 VDD P L=1.8e-07 W=6.85e-07 $X=1225 $Y=2555 $D=16
M6 10 A2 ZN VDD P L=1.8e-07 W=6.85e-07 $X=1945 $Y=2555 $D=16
M7 VDD B1 10 VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2890 $D=16
.ENDS
***************************************
.SUBCKT XNR3D0BWP7T A2 A1 A3 VDD VSS ZN
** N=16 EP=6 IP=0 FDC=22
M0 VSS A2 7 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=845 $D=0
M1 13 8 VSS VSS N L=1.8e-07 W=5e-07 $X=1500 $Y=845 $D=0
M2 9 7 13 VSS N L=1.8e-07 W=5e-07 $X=2045 $Y=845 $D=0
M3 8 A2 9 VSS N L=1.8e-07 W=5e-07 $X=2825 $Y=845 $D=0
M4 VSS A1 8 VSS N L=1.8e-07 W=7.05e-07 $X=3545 $Y=640 $D=0
M5 VSS 9 10 VSS N L=1.8e-07 W=5e-07 $X=5115 $Y=460 $D=0
M6 14 11 VSS VSS N L=1.8e-07 W=5e-07 $X=5915 $Y=845 $D=0
M7 12 10 14 VSS N L=1.8e-07 W=5e-07 $X=6345 $Y=845 $D=0
M8 11 9 12 VSS N L=1.8e-07 W=5e-07 $X=7205 $Y=440 $D=0
M9 VSS A3 11 VSS N L=1.8e-07 W=5e-07 $X=7965 $Y=440 $D=0
M10 ZN 12 VSS VSS N L=1.8e-07 W=5e-07 $X=8720 $Y=440 $D=0
M11 VDD A2 7 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2645 $D=16
M12 15 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1420 $Y=2435 $D=16
M13 9 A2 15 VDD P L=1.8e-07 W=6.85e-07 $X=1900 $Y=2435 $D=16
M14 8 7 9 VDD P L=1.8e-07 W=6.85e-07 $X=2745 $Y=2435 $D=16
M15 VDD A1 8 VDD P L=1.8e-07 W=6.85e-07 $X=3545 $Y=2435 $D=16
M16 VDD 9 10 VDD P L=1.8e-07 W=6.85e-07 $X=5115 $Y=2815 $D=16
M17 16 11 VDD VDD P L=1.8e-07 W=6.85e-07 $X=5915 $Y=2445 $D=16
M18 12 9 16 VDD P L=1.8e-07 W=6.85e-07 $X=6425 $Y=2445 $D=16
M19 11 10 12 VDD P L=1.8e-07 W=6.85e-07 $X=7145 $Y=2445 $D=16
M20 VDD A3 11 VDD P L=1.8e-07 W=6.85e-07 $X=7905 $Y=2205 $D=16
M21 ZN 12 VDD VDD P L=1.8e-07 W=6.85e-07 $X=8720 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKBD0BWP7T I VSS VDD Z
** N=5 EP=4 IP=0 FDC=4
M0 VSS I 5 VSS N L=1.8e-07 W=4.2e-07 $X=620 $Y=445 $D=0
M1 Z 5 VSS VSS N L=1.8e-07 W=4.2e-07 $X=1440 $Y=445 $D=0
M2 VDD I 5 VDD P L=1.8e-07 W=1.27e-06 $X=620 $Y=2290 $D=16
M3 Z 5 VDD VDD P L=1.8e-07 W=1.13e-06 $X=1440 $Y=2430 $D=16
.ENDS
***************************************
.SUBCKT AO211D1BWP7T A1 A2 B C VDD VSS Z
** N=11 EP=7 IP=0 FDC=10
M0 10 A1 9 VSS N L=1.8e-07 W=1e-06 $X=660 $Y=345 $D=0
M1 VSS A2 10 VSS N L=1.8e-07 W=1e-06 $X=1140 $Y=345 $D=0
M2 9 B VSS VSS N L=1.8e-07 W=1e-06 $X=2100 $Y=345 $D=0
M3 VSS C 9 VSS N L=1.8e-07 W=1e-06 $X=2830 $Y=345 $D=0
M4 Z 9 VSS VSS N L=1.8e-07 W=1e-06 $X=3595 $Y=345 $D=0
M5 9 A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M6 8 A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=1380 $Y=2205 $D=16
M7 11 B 8 VDD P L=1.8e-07 W=1.37e-06 $X=2100 $Y=2205 $D=16
M8 VDD C 11 VDD P L=1.8e-07 W=1.37e-06 $X=2805 $Y=2205 $D=16
M9 Z 9 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3595 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR2D1BWP7T A2 VDD ZN A1 VSS
** N=6 EP=5 IP=0 FDC=4
M0 ZN A2 VSS VSS N L=1.8e-07 W=1e-06 $X=660 $Y=345 $D=0
M1 VSS A1 ZN VSS N L=1.8e-07 W=1e-06 $X=1420 $Y=345 $D=0
M2 6 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M3 ZN A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=1260 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AOI21D0BWP7T A2 ZN A1 B VSS VDD
** N=8 EP=6 IP=0 FDC=6
M0 8 A2 VSS VSS N L=1.8e-07 W=5e-07 $X=630 $Y=460 $D=0
M1 ZN A1 8 VSS N L=1.8e-07 W=5e-07 $X=1250 $Y=460 $D=0
M2 VSS B ZN VSS N L=1.8e-07 W=5e-07 $X=1975 $Y=460 $D=0
M3 ZN A2 7 VDD P L=1.8e-07 W=6.85e-07 $X=630 $Y=2275 $D=16
M4 7 A1 ZN VDD P L=1.8e-07 W=6.85e-07 $X=1355 $Y=2275 $D=16
M5 VDD B 7 VDD P L=1.8e-07 W=6.85e-07 $X=2075 $Y=2275 $D=16
.ENDS
***************************************
.SUBCKT NR4D1BWP7T ZN A1 A2 A4 VDD VSS A3
** N=13 EP=7 IP=0 FDC=12
M0 ZN A1 VSS VSS N L=1.8e-07 W=1e-06 $X=1830 $Y=345 $D=0
M1 VSS A2 ZN VSS N L=1.8e-07 W=1e-06 $X=2550 $Y=345 $D=0
M2 ZN A3 VSS VSS N L=1.8e-07 W=1e-06 $X=3360 $Y=345 $D=0
M3 VSS A4 ZN VSS N L=1.8e-07 W=1e-06 $X=4080 $Y=345 $D=0
M4 9 A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M5 ZN A1 9 VDD P L=1.8e-07 W=1.37e-06 $X=1160 $Y=2205 $D=16
M6 10 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1880 $Y=2205 $D=16
M7 11 A2 10 VDD P L=1.8e-07 W=1.37e-06 $X=2470 $Y=2205 $D=16
M8 12 A3 11 VDD P L=1.8e-07 W=1.37e-06 $X=3060 $Y=2205 $D=16
M9 VDD A4 12 VDD P L=1.8e-07 W=1.37e-06 $X=3650 $Y=2205 $D=16
M10 13 A4 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4370 $Y=2205 $D=16
M11 8 A3 13 VDD P L=1.8e-07 W=1.37e-06 $X=4800 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AN3D1BWP7T A1 A2 A3 VDD VSS Z
** N=9 EP=6 IP=0 FDC=8
M0 8 A1 7 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=345 $D=0
M1 9 A2 8 VSS N L=1.8e-07 W=5e-07 $X=1205 $Y=345 $D=0
M2 VSS A3 9 VSS N L=1.8e-07 W=5e-07 $X=1790 $Y=345 $D=0
M3 Z 7 VSS VSS N L=1.8e-07 W=1e-06 $X=2560 $Y=345 $D=0
M4 VDD A1 7 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2205 $D=16
M5 7 A2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1230 $Y=2205 $D=16
M6 VDD A3 7 VDD P L=1.8e-07 W=6.85e-07 $X=1950 $Y=2205 $D=16
M7 Z 7 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2560 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AOI31D2BWP7T B VDD ZN A1 A2 A3 VSS
** N=12 EP=7 IP=0 FDC=16
M0 ZN B VSS VSS N L=1.8e-07 W=1e-06 $X=645 $Y=345 $D=0
M1 VSS B ZN VSS N L=1.8e-07 W=1e-06 $X=1370 $Y=345 $D=0
M2 9 A3 VSS VSS N L=1.8e-07 W=1e-06 $X=2490 $Y=345 $D=0
M3 10 A2 9 VSS N L=1.8e-07 W=8.45e-07 $X=3160 $Y=345 $D=0
M4 ZN A1 10 VSS N L=1.8e-07 W=8.45e-07 $X=3830 $Y=345 $D=0
M5 11 A1 ZN VSS N L=1.8e-07 W=8.8e-07 $X=4630 $Y=345 $D=0
M6 12 A2 11 VSS N L=1.8e-07 W=8.8e-07 $X=5230 $Y=345 $D=0
M7 VSS A3 12 VSS N L=1.8e-07 W=8.8e-07 $X=5830 $Y=345 $D=0
M8 VDD B 8 VDD P L=1.8e-07 W=1.3e-06 $X=645 $Y=2275 $D=16
M9 8 B VDD VDD P L=1.8e-07 W=1.3e-06 $X=1370 $Y=2275 $D=16
M10 ZN A3 8 VDD P L=1.8e-07 W=1.3e-06 $X=2090 $Y=2275 $D=16
M11 8 A3 ZN VDD P L=1.8e-07 W=1.3e-06 $X=2810 $Y=2275 $D=16
M12 ZN A1 8 VDD P L=1.8e-07 W=1.3e-06 $X=3610 $Y=2275 $D=16
M13 8 A1 ZN VDD P L=1.8e-07 W=1.3e-06 $X=4330 $Y=2275 $D=16
M14 ZN A2 8 VDD P L=1.8e-07 W=1.3e-06 $X=5150 $Y=2275 $D=16
M15 8 A2 ZN VDD P L=1.8e-07 W=1.3e-06 $X=5870 $Y=2275 $D=16
.ENDS
***************************************
.SUBCKT OR4D1BWP7T A4 A3 A2 A1 VDD VSS Z
** N=11 EP=7 IP=0 FDC=10
M0 8 A4 VSS VSS N L=1.8e-07 W=5e-07 $X=675 $Y=345 $D=0
M1 VSS A3 8 VSS N L=1.8e-07 W=5e-07 $X=1395 $Y=345 $D=0
M2 8 A2 VSS VSS N L=1.8e-07 W=5e-07 $X=2125 $Y=345 $D=0
M3 VSS A1 8 VSS N L=1.8e-07 W=5e-07 $X=2845 $Y=345 $D=0
M4 Z 8 VSS VSS N L=1.8e-07 W=1e-06 $X=3645 $Y=345 $D=0
M5 9 A4 8 VDD P L=1.8e-07 W=1.37e-06 $X=725 $Y=2205 $D=16
M6 10 A3 9 VDD P L=1.8e-07 W=1.37e-06 $X=1325 $Y=2205 $D=16
M7 11 A2 10 VDD P L=1.8e-07 W=1.37e-06 $X=1925 $Y=2205 $D=16
M8 VDD A1 11 VDD P L=1.8e-07 W=1.37e-06 $X=2525 $Y=2205 $D=16
M9 Z 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3275 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OA31D0BWP7T A1 A2 A3 B VSS VDD Z
** N=11 EP=7 IP=0 FDC=10
M0 8 A1 9 VSS N L=1.8e-07 W=5e-07 $X=665 $Y=750 $D=0
M1 9 A2 8 VSS N L=1.8e-07 W=5e-07 $X=1385 $Y=750 $D=0
M2 8 A3 9 VSS N L=1.8e-07 W=5e-07 $X=2165 $Y=750 $D=0
M3 VSS B 8 VSS N L=1.8e-07 W=5e-07 $X=2910 $Y=750 $D=0
M4 Z 9 VSS VSS N L=1.8e-07 W=5e-07 $X=3670 $Y=750 $D=0
M5 10 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=665 $Y=2860 $D=16
M6 11 A2 10 VDD P L=1.8e-07 W=6.85e-07 $X=1385 $Y=2860 $D=16
M7 9 A3 11 VDD P L=1.8e-07 W=6.85e-07 $X=2105 $Y=2860 $D=16
M8 VDD B 9 VDD P L=1.8e-07 W=6.85e-07 $X=2910 $Y=2860 $D=16
M9 Z 9 VDD VDD P L=1.8e-07 W=6.85e-07 $X=3670 $Y=2860 $D=16
.ENDS
***************************************
.SUBCKT AOI21D2BWP7T B VDD ZN A1 A2 VSS
** N=9 EP=6 IP=0 FDC=12
M0 ZN B VSS VSS N L=1.8e-07 W=1e-06 $X=625 $Y=345 $D=0
M1 VSS B ZN VSS N L=1.8e-07 W=1e-06 $X=1345 $Y=345 $D=0
M2 8 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=2145 $Y=345 $D=0
M3 ZN A1 8 VSS N L=1.8e-07 W=1e-06 $X=2800 $Y=345 $D=0
M4 9 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=3520 $Y=345 $D=0
M5 VSS A2 9 VSS N L=1.8e-07 W=1e-06 $X=4240 $Y=345 $D=0
M6 VDD B 7 VDD P L=1.8e-07 W=1.37e-06 $X=625 $Y=2205 $D=16
M7 7 B VDD VDD P L=1.8e-07 W=1.37e-06 $X=1345 $Y=2205 $D=16
M8 ZN A2 7 VDD P L=1.8e-07 W=1.37e-06 $X=2080 $Y=2205 $D=16
M9 7 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2800 $Y=2205 $D=16
M10 ZN A1 7 VDD P L=1.8e-07 W=1.37e-06 $X=3520 $Y=2205 $D=16
M11 7 A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4240 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ND2D1BWP7T A2 VSS ZN A1 VDD
** N=6 EP=5 IP=0 FDC=4
M0 6 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=660 $Y=345 $D=0
M1 ZN A1 6 VSS N L=1.8e-07 W=1e-06 $X=1300 $Y=345 $D=0
M2 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M3 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1380 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OAI211D1BWP7T C VSS B A1 VDD ZN A2
** N=10 EP=7 IP=0 FDC=8
M0 9 C VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 8 B 9 VSS N L=1.8e-07 W=1e-06 $X=1120 $Y=345 $D=0
M2 ZN A1 8 VSS N L=1.8e-07 W=1e-06 $X=1840 $Y=345 $D=0
M3 8 A2 ZN VSS N L=1.8e-07 W=1e-06 $X=2560 $Y=345 $D=0
M4 ZN C VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M5 VDD B ZN VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M6 10 A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M7 ZN A2 10 VDD P L=1.8e-07 W=1.37e-06 $X=2560 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR4D2BWP7T A4 VDD A3 A2 A1 VSS ZN
** N=10 EP=7 IP=0 FDC=32
M0 VSS A4 ZN VSS N L=1.8e-07 W=5e-07 $X=620 $Y=345 $D=0
M1 ZN A4 VSS VSS N L=1.8e-07 W=5e-07 $X=1340 $Y=345 $D=0
M2 VSS A4 ZN VSS N L=1.8e-07 W=5e-07 $X=2060 $Y=345 $D=0
M3 ZN A4 VSS VSS N L=1.8e-07 W=5e-07 $X=2780 $Y=345 $D=0
M4 VSS A3 ZN VSS N L=1.8e-07 W=5e-07 $X=3500 $Y=345 $D=0
M5 ZN A3 VSS VSS N L=1.8e-07 W=5e-07 $X=4220 $Y=345 $D=0
M6 VSS A3 ZN VSS N L=1.8e-07 W=5e-07 $X=4940 $Y=345 $D=0
M7 ZN A3 VSS VSS N L=1.8e-07 W=5e-07 $X=5660 $Y=345 $D=0
M8 VSS A2 ZN VSS N L=1.8e-07 W=5e-07 $X=7040 $Y=345 $D=0
M9 ZN A2 VSS VSS N L=1.8e-07 W=5e-07 $X=7760 $Y=345 $D=0
M10 VSS A2 ZN VSS N L=1.8e-07 W=5e-07 $X=8480 $Y=345 $D=0
M11 ZN A2 VSS VSS N L=1.8e-07 W=5e-07 $X=9200 $Y=345 $D=0
M12 VSS A1 ZN VSS N L=1.8e-07 W=5e-07 $X=9920 $Y=345 $D=0
M13 ZN A1 VSS VSS N L=1.8e-07 W=5e-07 $X=10640 $Y=345 $D=0
M14 VSS A1 ZN VSS N L=1.8e-07 W=5e-07 $X=11360 $Y=345 $D=0
M15 ZN A1 VSS VSS N L=1.8e-07 W=5e-07 $X=12080 $Y=345 $D=0
M16 VDD A4 8 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M17 8 A4 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M18 VDD A4 8 VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M19 8 A4 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M20 9 A3 8 VDD P L=1.8e-07 W=1.37e-06 $X=3500 $Y=2205 $D=16
M21 8 A3 9 VDD P L=1.8e-07 W=1.37e-06 $X=4220 $Y=2205 $D=16
M22 9 A3 8 VDD P L=1.8e-07 W=1.37e-06 $X=4940 $Y=2205 $D=16
M23 8 A3 9 VDD P L=1.8e-07 W=1.37e-06 $X=5660 $Y=2205 $D=16
M24 9 A2 10 VDD P L=1.8e-07 W=1.37e-06 $X=7040 $Y=2205 $D=16
M25 10 A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=7760 $Y=2205 $D=16
M26 9 A2 10 VDD P L=1.8e-07 W=1.37e-06 $X=8480 $Y=2205 $D=16
M27 10 A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=9200 $Y=2205 $D=16
M28 ZN A1 10 VDD P L=1.8e-07 W=1.37e-06 $X=9920 $Y=2205 $D=16
M29 10 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=10640 $Y=2205 $D=16
M30 ZN A1 10 VDD P L=1.8e-07 W=1.37e-06 $X=11360 $Y=2205 $D=16
M31 10 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=12080 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR2XD0BWP7T A2 VDD A1 ZN VSS
** N=6 EP=5 IP=0 FDC=4
M0 ZN A2 VSS VSS N L=1.8e-07 W=5e-07 $X=720 $Y=360 $D=0
M1 VSS A1 ZN VSS N L=1.8e-07 W=5e-07 $X=1440 $Y=360 $D=0
M2 6 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=720 $Y=2205 $D=16
M3 ZN A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=1320 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OA22D0BWP7T B2 B1 A1 A2 VDD VSS Z
** N=11 EP=7 IP=0 FDC=10
M0 9 B2 VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=805 $D=0
M1 8 A1 9 VSS N L=1.8e-07 W=5e-07 $X=1360 $Y=805 $D=0
M2 9 A2 8 VSS N L=1.8e-07 W=5e-07 $X=2240 $Y=805 $D=0
M3 VSS B1 9 VSS N L=1.8e-07 W=5e-07 $X=2960 $Y=805 $D=0
M4 Z 8 VSS VSS N L=1.8e-07 W=5e-07 $X=3680 $Y=805 $D=0
M5 10 B2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2890 $D=16
M6 8 B1 10 VDD P L=1.8e-07 W=6.85e-07 $X=1180 $Y=2890 $D=16
M7 11 A1 8 VDD P L=1.8e-07 W=6.85e-07 $X=1900 $Y=2890 $D=16
M8 VDD A2 11 VDD P L=1.8e-07 W=6.85e-07 $X=2520 $Y=2890 $D=16
M9 Z 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=3630 $Y=2890 $D=16
.ENDS
***************************************
.SUBCKT ND4D1BWP7T A4 VSS A3 A2 A1 ZN VDD
** N=10 EP=7 IP=0 FDC=8
M0 8 A4 VSS VSS N L=1.8e-07 W=1e-06 $X=660 $Y=345 $D=0
M1 9 A3 8 VSS N L=1.8e-07 W=1e-06 $X=1300 $Y=345 $D=0
M2 10 A2 9 VSS N L=1.8e-07 W=1e-06 $X=1940 $Y=345 $D=0
M3 ZN A1 10 VSS N L=1.8e-07 W=1e-06 $X=2580 $Y=345 $D=0
M4 ZN A4 VDD VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M5 VDD A3 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1380 $Y=2205 $D=16
M6 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2100 $Y=2205 $D=16
M7 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2820 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OAI31D1BWP7T A1 A2 ZN A3 B VSS VDD
** N=10 EP=7 IP=0 FDC=8
M0 8 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=680 $Y=345 $D=0
M1 ZN A2 8 VSS N L=1.8e-07 W=1e-06 $X=1400 $Y=345 $D=0
M2 8 A3 ZN VSS N L=1.8e-07 W=1e-06 $X=2160 $Y=345 $D=0
M3 VSS B 8 VSS N L=1.8e-07 W=1e-06 $X=2930 $Y=345 $D=0
M4 9 A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=680 $Y=2205 $D=16
M5 10 A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=1400 $Y=2205 $D=16
M6 ZN A3 10 VDD P L=1.8e-07 W=1.37e-06 $X=2120 $Y=2205 $D=16
M7 VDD B ZN VDD P L=1.8e-07 W=1.37e-06 $X=2930 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AOI31D0BWP7T A3 A2 A1 ZN B VSS VDD
** N=10 EP=7 IP=0 FDC=8
M0 8 A3 VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=480 $D=0
M1 9 A2 8 VSS N L=1.8e-07 W=5e-07 $X=1210 $Y=480 $D=0
M2 ZN A1 9 VSS N L=1.8e-07 W=5e-07 $X=1800 $Y=480 $D=0
M3 VSS B ZN VSS N L=1.8e-07 W=5e-07 $X=2560 $Y=480 $D=0
M4 10 A3 ZN VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2250 $D=16
M5 ZN A2 10 VDD P L=1.8e-07 W=6.85e-07 $X=1220 $Y=2250 $D=16
M6 10 A1 ZN VDD P L=1.8e-07 W=6.85e-07 $X=1945 $Y=2250 $D=16
M7 VDD B 10 VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2250 $D=16
.ENDS
***************************************
.SUBCKT ND3D0BWP7T A3 VSS A2 A1 VDD ZN
** N=8 EP=6 IP=0 FDC=6
M0 7 A3 VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=500 $D=0
M1 8 A2 7 VSS N L=1.8e-07 W=5e-07 $X=1245 $Y=500 $D=0
M2 ZN A1 8 VSS N L=1.8e-07 W=5e-07 $X=1870 $Y=500 $D=0
M3 ZN A3 VDD VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2735 $D=16
M4 VDD A2 ZN VDD P L=1.8e-07 W=6.85e-07 $X=1340 $Y=2735 $D=16
M5 ZN A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=2000 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR4D0BWP7T A4 VSS VDD A3 A2 ZN A1
** N=10 EP=7 IP=0 FDC=8
M0 ZN A4 VSS VSS N L=1.8e-07 W=5e-07 $X=625 $Y=725 $D=0
M1 VSS A3 ZN VSS N L=1.8e-07 W=5e-07 $X=1345 $Y=725 $D=0
M2 ZN A2 VSS VSS N L=1.8e-07 W=5e-07 $X=1945 $Y=725 $D=0
M3 VSS A1 ZN VSS N L=1.8e-07 W=5e-07 $X=2680 $Y=725 $D=0
M4 8 A4 VDD VDD P L=1.8e-07 W=1.37e-06 $X=625 $Y=2205 $D=16
M5 9 A3 8 VDD P L=1.8e-07 W=1.37e-06 $X=1265 $Y=2205 $D=16
M6 10 A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=1905 $Y=2205 $D=16
M7 ZN A1 10 VDD P L=1.8e-07 W=1.37e-06 $X=2545 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR2D2BWP7T A2 A1 VDD ZN VSS
** N=6 EP=5 IP=0 FDC=8
M0 ZN A2 VSS VSS N L=1.8e-07 W=1e-06 $X=660 $Y=345 $D=0
M1 VSS A2 ZN VSS N L=1.8e-07 W=1e-06 $X=1380 $Y=345 $D=0
M2 ZN A1 VSS VSS N L=1.8e-07 W=1e-06 $X=2240 $Y=345 $D=0
M3 VSS A1 ZN VSS N L=1.8e-07 W=1e-06 $X=2960 $Y=345 $D=0
M4 VDD A2 6 VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M5 6 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1380 $Y=2205 $D=16
M6 ZN A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=2240 $Y=2205 $D=16
M7 6 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2960 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AN4D1BWP7T A1 A2 A3 A4 VDD VSS Z
** N=11 EP=7 IP=0 FDC=10
M0 9 A1 8 VSS N L=1.8e-07 W=5e-07 $X=625 $Y=345 $D=0
M1 10 A2 9 VSS N L=1.8e-07 W=5e-07 $X=1205 $Y=345 $D=0
M2 11 A3 10 VSS N L=1.8e-07 W=5e-07 $X=1785 $Y=345 $D=0
M3 VSS A4 11 VSS N L=1.8e-07 W=5e-07 $X=2365 $Y=345 $D=0
M4 Z 8 VSS VSS N L=1.8e-07 W=1e-06 $X=3105 $Y=345 $D=0
M5 8 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=460 $Y=2205 $D=16
M6 VDD A2 8 VDD P L=1.8e-07 W=6.85e-07 $X=1185 $Y=2205 $D=16
M7 8 A3 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1785 $Y=2205 $D=16
M8 VDD A4 8 VDD P L=1.8e-07 W=6.85e-07 $X=2515 $Y=2205 $D=16
M9 Z 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3115 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT BUFFD0BWP7T I VSS VDD Z
** N=5 EP=4 IP=0 FDC=4
M0 VSS I 5 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=555 $D=0
M1 Z 5 VSS VSS N L=1.8e-07 W=5e-07 $X=1420 $Y=555 $D=0
M2 VDD I 5 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2850 $D=16
M3 Z 5 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1420 $Y=2850 $D=16
.ENDS
***************************************
.SUBCKT AOI31D1BWP7T A3 A2 ZN A1 B VDD VSS
** N=10 EP=7 IP=0 FDC=8
M0 9 A3 VSS VSS N L=1.8e-07 W=1e-06 $X=680 $Y=345 $D=0
M1 10 A2 9 VSS N L=1.8e-07 W=1e-06 $X=1385 $Y=345 $D=0
M2 ZN A1 10 VSS N L=1.8e-07 W=1e-06 $X=2090 $Y=345 $D=0
M3 VSS B ZN VSS N L=1.8e-07 W=1e-06 $X=2930 $Y=345 $D=0
M4 8 A3 ZN VDD P L=1.8e-07 W=1.37e-06 $X=680 $Y=2205 $D=16
M5 ZN A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=1400 $Y=2205 $D=16
M6 8 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2160 $Y=2205 $D=16
M7 VDD B 8 VDD P L=1.8e-07 W=1.37e-06 $X=2930 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ND4D0BWP7T A4 VSS A3 A2 A1 ZN VDD
** N=10 EP=7 IP=0 FDC=8
M0 8 A4 VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=360 $D=0
M1 9 A3 8 VSS N L=1.8e-07 W=5e-07 $X=1240 $Y=360 $D=0
M2 10 A2 9 VSS N L=1.8e-07 W=5e-07 $X=1860 $Y=360 $D=0
M3 ZN A1 10 VSS N L=1.8e-07 W=5e-07 $X=2480 $Y=360 $D=0
M4 ZN A4 VDD VDD P L=1.8e-07 W=6.85e-07 $X=575 $Y=2235 $D=16
M5 VDD A3 ZN VDD P L=1.8e-07 W=6.85e-07 $X=1295 $Y=2235 $D=16
M6 ZN A2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1955 $Y=2235 $D=16
M7 VDD A1 ZN VDD P L=1.8e-07 W=6.85e-07 $X=2690 $Y=2235 $D=16
.ENDS
***************************************
.SUBCKT IND3D1BWP7T A1 VSS B1 VDD B2 ZN
** N=9 EP=6 IP=0 FDC=8
M0 VSS A1 7 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=360 $D=0
M1 8 7 VSS VSS N L=1.8e-07 W=1e-06 $X=1420 $Y=345 $D=0
M2 9 B1 8 VSS N L=1.8e-07 W=1e-06 $X=1980 $Y=345 $D=0
M3 ZN B2 9 VSS N L=1.8e-07 W=1e-06 $X=2540 $Y=345 $D=0
M4 VDD A1 7 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2205 $D=16
M5 ZN 7 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1225 $Y=2205 $D=16
M6 VDD B1 ZN VDD P L=1.8e-07 W=8.35e-07 $X=1945 $Y=2205 $D=16
M7 ZN B2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2560 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR2D1P5BWP7T A1 ZN A2 VDD VSS
** N=7 EP=5 IP=0 FDC=8
M0 ZN A2 VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS A1 ZN VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 ZN A1 VSS VSS N L=1.8e-07 W=5e-07 $X=2080 $Y=345 $D=0
M3 VSS A2 ZN VSS N L=1.8e-07 W=5e-07 $X=2800 $Y=345 $D=0
M4 6 A2 VDD VDD P L=1.8e-07 W=1.03e-06 $X=620 $Y=2545 $D=16
M5 ZN A1 6 VDD P L=1.8e-07 W=1.03e-06 $X=1220 $Y=2545 $D=16
M6 7 A1 ZN VDD P L=1.8e-07 W=1.03e-06 $X=1940 $Y=2545 $D=16
M7 VDD A2 7 VDD P L=1.8e-07 W=1.03e-06 $X=2800 $Y=2545 $D=16
.ENDS
***************************************
.SUBCKT OA21D0BWP7T A2 A1 B VDD VSS Z
** N=9 EP=6 IP=0 FDC=8
M0 7 A2 8 VSS N L=1.8e-07 W=5e-07 $X=460 $Y=750 $D=0
M1 8 A1 7 VSS N L=1.8e-07 W=5e-07 $X=1180 $Y=750 $D=0
M2 VSS B 8 VSS N L=1.8e-07 W=5e-07 $X=1840 $Y=455 $D=0
M3 Z 7 VSS VSS N L=1.8e-07 W=5e-07 $X=2560 $Y=455 $D=0
M4 9 A2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=460 $Y=2350 $D=16
M5 7 A1 9 VDD P L=1.8e-07 W=6.85e-07 $X=1120 $Y=2350 $D=16
M6 VDD B 7 VDD P L=1.8e-07 W=6.85e-07 $X=1840 $Y=2350 $D=16
M7 Z 7 VDD VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2585 $D=16
.ENDS
***************************************
.SUBCKT INR4D0BWP7T A1 VDD B1 B2 B3 ZN VSS
** N=11 EP=7 IP=0 FDC=10
M0 VSS A1 8 VSS N L=1.8e-07 W=4.2e-07 $X=620 $Y=425 $D=0
M1 ZN 8 VSS VSS N L=1.8e-07 W=5e-07 $X=1340 $Y=345 $D=0
M2 VSS B1 ZN VSS N L=1.8e-07 W=5e-07 $X=2160 $Y=345 $D=0
M3 ZN B2 VSS VSS N L=1.8e-07 W=5e-07 $X=2960 $Y=345 $D=0
M4 VSS B3 ZN VSS N L=1.8e-07 W=5e-07 $X=3680 $Y=345 $D=0
M5 VDD A1 8 VDD P L=1.8e-07 W=4.2e-07 $X=620 $Y=2470 $D=16
M6 9 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1440 $Y=2205 $D=16
M7 10 B1 9 VDD P L=1.8e-07 W=1.37e-06 $X=2160 $Y=2205 $D=16
M8 11 B2 10 VDD P L=1.8e-07 W=1.37e-06 $X=2880 $Y=2205 $D=16
M9 ZN B3 11 VDD P L=1.8e-07 W=1.37e-06 $X=3600 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IND3D0BWP7T A1 VSS B1 B2 VDD ZN
** N=9 EP=6 IP=0 FDC=8
M0 VSS A1 7 VSS N L=1.8e-07 W=4.2e-07 $X=620 $Y=460 $D=0
M1 8 7 VSS VSS N L=1.8e-07 W=5e-07 $X=1340 $Y=460 $D=0
M2 9 B1 8 VSS N L=1.8e-07 W=5e-07 $X=1940 $Y=460 $D=0
M3 ZN B2 9 VSS N L=1.8e-07 W=5e-07 $X=2540 $Y=460 $D=0
M4 VDD A1 7 VDD P L=1.8e-07 W=4.2e-07 $X=620 $Y=2890 $D=16
M5 ZN 7 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1225 $Y=2320 $D=16
M6 VDD B1 ZN VDD P L=1.8e-07 W=6.85e-07 $X=1945 $Y=2320 $D=16
M7 ZN B2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2320 $D=16
.ENDS
***************************************
.SUBCKT NR3D1BWP7T A1 VSS A2 A3 ZN VDD
** N=10 EP=6 IP=0 FDC=9
M0 ZN A3 VSS VSS N L=1.8e-07 W=1e-06 $X=640 $Y=345 $D=0
M1 VSS A2 ZN VSS N L=1.8e-07 W=1e-06 $X=1360 $Y=345 $D=0
M2 ZN A1 VSS VSS N L=1.8e-07 W=1e-06 $X=2160 $Y=345 $D=0
M3 7 A3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=640 $Y=2205 $D=16
M4 8 A2 7 VDD P L=1.8e-07 W=1.37e-06 $X=1230 $Y=2205 $D=16
M5 ZN A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=1820 $Y=2205 $D=16
M6 9 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2540 $Y=2205 $D=16
M7 10 A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=3095 $Y=2205 $D=16
M8 VDD A3 10 VDD P L=1.8e-07 W=1.37e-06 $X=3650 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IND4D0BWP7T A1 VSS B1 B2 ZN B3 VDD
** N=11 EP=7 IP=0 FDC=10
M0 VSS A1 8 VSS N L=1.8e-07 W=4.2e-07 $X=620 $Y=425 $D=0
M1 9 8 VSS VSS N L=1.8e-07 W=5e-07 $X=1340 $Y=345 $D=0
M2 10 B1 9 VSS N L=1.8e-07 W=5e-07 $X=1930 $Y=345 $D=0
M3 11 B2 10 VSS N L=1.8e-07 W=5e-07 $X=2520 $Y=345 $D=0
M4 ZN B3 11 VSS N L=1.8e-07 W=5e-07 $X=3110 $Y=345 $D=0
M5 VDD A1 8 VDD P L=1.8e-07 W=4.2e-07 $X=620 $Y=2845 $D=16
M6 ZN 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1220 $Y=2320 $D=16
M7 VDD B1 ZN VDD P L=1.8e-07 W=6.85e-07 $X=1940 $Y=2320 $D=16
M8 ZN B2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=2540 $Y=2320 $D=16
M9 VDD B3 ZN VDD P L=1.8e-07 W=6.85e-07 $X=3260 $Y=2320 $D=16
.ENDS
***************************************
.SUBCKT IND4D1BWP7T A1 VSS B1 B2 ZN B3 VDD
** N=11 EP=7 IP=0 FDC=10
M0 VSS A1 8 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=500 $D=0
M1 9 8 VSS VSS N L=1.8e-07 W=1e-06 $X=1420 $Y=345 $D=0
M2 10 B1 9 VSS N L=1.8e-07 W=1e-06 $X=2140 $Y=345 $D=0
M3 11 B2 10 VSS N L=1.8e-07 W=1e-06 $X=2860 $Y=345 $D=0
M4 ZN B3 11 VSS N L=1.8e-07 W=1e-06 $X=3580 $Y=345 $D=0
M5 VDD A1 8 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2205 $D=16
M6 ZN 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1420 $Y=2205 $D=16
M7 VDD B1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2140 $Y=2205 $D=16
M8 ZN B2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2860 $Y=2205 $D=16
M9 VDD B3 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3580 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR4D3BWP7T A4 VDD A3 A2 A1 VSS ZN
** N=10 EP=7 IP=0 FDC=40
M0 VSS A4 ZN VSS N L=1.8e-07 W=6e-07 $X=830 $Y=345 $D=0
M1 ZN A4 VSS VSS N L=1.8e-07 W=6e-07 $X=1550 $Y=345 $D=0
M2 VSS A4 ZN VSS N L=1.8e-07 W=6e-07 $X=2270 $Y=345 $D=0
M3 ZN A4 VSS VSS N L=1.8e-07 W=6e-07 $X=2990 $Y=345 $D=0
M4 VSS A4 ZN VSS N L=1.8e-07 W=6e-07 $X=3710 $Y=345 $D=0
M5 ZN A3 VSS VSS N L=1.8e-07 W=6e-07 $X=4430 $Y=345 $D=0
M6 VSS A3 ZN VSS N L=1.8e-07 W=6e-07 $X=5150 $Y=345 $D=0
M7 ZN A3 VSS VSS N L=1.8e-07 W=6e-07 $X=5870 $Y=345 $D=0
M8 VSS A3 ZN VSS N L=1.8e-07 W=6e-07 $X=6590 $Y=345 $D=0
M9 ZN A3 VSS VSS N L=1.8e-07 W=6e-07 $X=7310 $Y=345 $D=0
M10 VSS A2 ZN VSS N L=1.8e-07 W=6e-07 $X=8030 $Y=345 $D=0
M11 ZN A2 VSS VSS N L=1.8e-07 W=6e-07 $X=8750 $Y=345 $D=0
M12 VSS A2 ZN VSS N L=1.8e-07 W=6e-07 $X=9470 $Y=345 $D=0
M13 ZN A2 VSS VSS N L=1.8e-07 W=6e-07 $X=10190 $Y=345 $D=0
M14 VSS A2 ZN VSS N L=1.8e-07 W=6e-07 $X=10910 $Y=345 $D=0
M15 ZN A1 VSS VSS N L=1.8e-07 W=6e-07 $X=11630 $Y=345 $D=0
M16 VSS A1 ZN VSS N L=1.8e-07 W=6e-07 $X=12350 $Y=345 $D=0
M17 ZN A1 VSS VSS N L=1.8e-07 W=6e-07 $X=13070 $Y=345 $D=0
M18 VSS A1 ZN VSS N L=1.8e-07 W=6e-07 $X=13790 $Y=345 $D=0
M19 ZN A1 VSS VSS N L=1.8e-07 W=6e-07 $X=14510 $Y=345 $D=0
M20 8 A4 VDD VDD P L=1.8e-07 W=1.34e-06 $X=830 $Y=2235 $D=16
M21 VDD A4 8 VDD P L=1.8e-07 W=1.72e-06 $X=1550 $Y=1855 $D=16
M22 8 A4 VDD VDD P L=1.8e-07 W=1.72e-06 $X=2270 $Y=1855 $D=16
M23 VDD A4 8 VDD P L=1.8e-07 W=1.72e-06 $X=2990 $Y=1855 $D=16
M24 8 A4 VDD VDD P L=1.8e-07 W=1.72e-06 $X=3710 $Y=1855 $D=16
M25 10 A3 8 VDD P L=1.8e-07 W=1.645e-06 $X=4430 $Y=1930 $D=16
M26 8 A3 10 VDD P L=1.8e-07 W=1.645e-06 $X=5150 $Y=1930 $D=16
M27 10 A3 8 VDD P L=1.8e-07 W=1.645e-06 $X=5870 $Y=1930 $D=16
M28 8 A3 10 VDD P L=1.8e-07 W=1.645e-06 $X=6590 $Y=1930 $D=16
M29 10 A3 8 VDD P L=1.8e-07 W=1.645e-06 $X=7310 $Y=1930 $D=16
M30 9 A2 10 VDD P L=1.8e-07 W=1.645e-06 $X=8030 $Y=1930 $D=16
M31 10 A2 9 VDD P L=1.8e-07 W=1.645e-06 $X=8750 $Y=1930 $D=16
M32 9 A2 10 VDD P L=1.8e-07 W=1.645e-06 $X=9470 $Y=1930 $D=16
M33 10 A2 9 VDD P L=1.8e-07 W=1.645e-06 $X=10190 $Y=1930 $D=16
M34 9 A2 10 VDD P L=1.8e-07 W=1.645e-06 $X=10910 $Y=1930 $D=16
M35 ZN A1 9 VDD P L=1.8e-07 W=1.72e-06 $X=11630 $Y=1855 $D=16
M36 9 A1 ZN VDD P L=1.8e-07 W=1.72e-06 $X=12350 $Y=1855 $D=16
M37 ZN A1 9 VDD P L=1.8e-07 W=1.72e-06 $X=13070 $Y=1855 $D=16
M38 9 A1 ZN VDD P L=1.8e-07 W=1.72e-06 $X=13790 $Y=1855 $D=16
M39 ZN A1 9 VDD P L=1.8e-07 W=1.34e-06 $X=14510 $Y=2235 $D=16
.ENDS
***************************************
.SUBCKT OR4D0BWP7T A4 A3 A2 A1 VDD VSS Z
** N=11 EP=7 IP=0 FDC=10
M0 8 A4 VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=480 $D=0
M1 VSS A3 8 VSS N L=1.8e-07 W=5e-07 $X=1340 $Y=480 $D=0
M2 8 A2 VSS VSS N L=1.8e-07 W=5e-07 $X=2140 $Y=480 $D=0
M3 VSS A1 8 VSS N L=1.8e-07 W=5e-07 $X=2860 $Y=480 $D=0
M4 Z 8 VSS VSS N L=1.8e-07 W=5e-07 $X=3660 $Y=480 $D=0
M5 9 A4 8 VDD P L=1.8e-07 W=6.85e-07 $X=725 $Y=2875 $D=16
M6 10 A3 9 VDD P L=1.8e-07 W=6.85e-07 $X=1325 $Y=2875 $D=16
M7 11 A2 10 VDD P L=1.8e-07 W=6.85e-07 $X=1925 $Y=2875 $D=16
M8 VDD A1 11 VDD P L=1.8e-07 W=6.85e-07 $X=2525 $Y=2875 $D=16
M9 Z 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=3660 $Y=2875 $D=16
.ENDS
***************************************
.SUBCKT INR4D1BWP7T B2 B1 B3 ZN A1 VSS VDD
** N=14 EP=7 IP=0 FDC=14
M0 ZN B1 VSS VSS N L=1.8e-07 W=7e-07 $X=620 $Y=345 $D=0
M1 VSS B2 ZN VSS N L=1.8e-07 W=7e-07 $X=1340 $Y=345 $D=0
M2 ZN 9 VSS VSS N L=1.8e-07 W=7e-07 $X=3230 $Y=345 $D=0
M3 VSS B3 ZN VSS N L=1.8e-07 W=7e-07 $X=3950 $Y=345 $D=0
M4 VSS A1 9 VSS N L=1.8e-07 W=5e-07 $X=5675 $Y=460 $D=0
M5 10 B1 8 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M6 VDD B2 10 VDD P L=1.8e-07 W=1.37e-06 $X=1100 $Y=2205 $D=16
M7 11 B2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1840 $Y=2205 $D=16
M8 12 B1 11 VDD P L=1.8e-07 W=1.37e-06 $X=2370 $Y=2205 $D=16
M9 13 9 12 VDD P L=1.8e-07 W=1.37e-06 $X=2900 $Y=2205 $D=16
M10 ZN B3 13 VDD P L=1.8e-07 W=1.37e-06 $X=3430 $Y=2205 $D=16
M11 14 B3 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4150 $Y=2205 $D=16
M12 8 9 14 VDD P L=1.8e-07 W=1.37e-06 $X=4580 $Y=2205 $D=16
M13 VDD A1 9 VDD P L=1.8e-07 W=6.85e-07 $X=5920 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INR3D1BWP7T A1 B2 VSS B1 ZN VDD
** N=11 EP=6 IP=0 FDC=11
M0 VSS A1 7 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 ZN 7 VSS VSS N L=1.8e-07 W=1e-06 $X=1390 $Y=345 $D=0
M2 VSS B1 ZN VSS N L=1.8e-07 W=1e-06 $X=2110 $Y=345 $D=0
M3 ZN B2 VSS VSS N L=1.8e-07 W=1e-06 $X=2910 $Y=345 $D=0
M4 VDD A1 7 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M5 8 7 VDD VDD P L=1.8e-07 W=1.245e-06 $X=1390 $Y=2330 $D=16
M6 9 B1 8 VDD P L=1.8e-07 W=1.245e-06 $X=1940 $Y=2330 $D=16
M7 ZN B2 9 VDD P L=1.8e-07 W=1.245e-06 $X=2490 $Y=2330 $D=16
M8 10 B2 ZN VDD P L=1.8e-07 W=1.245e-06 $X=3230 $Y=2330 $D=16
M9 11 B1 10 VDD P L=1.8e-07 W=1.245e-06 $X=3735 $Y=2330 $D=16
M10 VDD 7 11 VDD P L=1.8e-07 W=1.245e-06 $X=4240 $Y=2330 $D=16
.ENDS
***************************************
.SUBCKT INR2D2BWP7T A1 B1 ZN VDD VSS
** N=8 EP=5 IP=0 FDC=10
M0 VSS A1 6 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 ZN 6 VSS VSS N L=1.8e-07 W=1e-06 $X=1480 $Y=345 $D=0
M2 VSS B1 ZN VSS N L=1.8e-07 W=1e-06 $X=2200 $Y=345 $D=0
M3 ZN B1 VSS VSS N L=1.8e-07 W=1e-06 $X=2960 $Y=345 $D=0
M4 VSS 6 ZN VSS N L=1.8e-07 W=1e-06 $X=3680 $Y=345 $D=0
M5 VDD A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M6 7 6 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1480 $Y=2205 $D=16
M7 ZN B1 7 VDD P L=1.8e-07 W=1.37e-06 $X=2200 $Y=2205 $D=16
M8 8 B1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2960 $Y=2205 $D=16
M9 VDD 6 8 VDD P L=1.8e-07 W=1.37e-06 $X=3680 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR2XD1BWP7T A2 VDD ZN VSS A1
** N=6 EP=5 IP=0 FDC=6
M0 ZN A2 VSS VSS N L=1.8e-07 W=1e-06 $X=1600 $Y=345 $D=0
M1 VSS A1 ZN VSS N L=1.8e-07 W=1e-06 $X=2320 $Y=345 $D=0
M2 VDD A2 6 VDD P L=1.8e-07 W=1.37e-06 $X=880 $Y=2205 $D=16
M3 6 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1600 $Y=2205 $D=16
M4 ZN A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=2320 $Y=2205 $D=16
M5 6 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3040 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IND2D1BWP7T A1 VSS ZN B1 VDD
** N=7 EP=5 IP=0 FDC=6
M0 VSS A1 6 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=565 $D=0
M1 7 6 VSS VSS N L=1.8e-07 W=1e-06 $X=1420 $Y=345 $D=0
M2 ZN B1 7 VSS N L=1.8e-07 W=1e-06 $X=2000 $Y=345 $D=0
M3 VDD A1 6 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2205 $D=16
M4 ZN 6 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1280 $Y=2205 $D=16
M5 VDD B1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2000 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OR4XD1BWP7T A4 A3 A2 A1 VDD VSS Z
** N=11 EP=7 IP=0 FDC=10
M0 8 A4 VSS VSS N L=1.8e-07 W=1e-06 $X=660 $Y=345 $D=0
M1 VSS A3 8 VSS N L=1.8e-07 W=1e-06 $X=1395 $Y=345 $D=0
M2 8 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=2115 $Y=345 $D=0
M3 VSS A1 8 VSS N L=1.8e-07 W=1e-06 $X=2835 $Y=345 $D=0
M4 Z 8 VSS VSS N L=1.8e-07 W=1e-06 $X=3555 $Y=345 $D=0
M5 9 A4 8 VDD P L=1.8e-07 W=1.37e-06 $X=705 $Y=2205 $D=16
M6 10 A3 9 VDD P L=1.8e-07 W=1.37e-06 $X=1335 $Y=2205 $D=16
M7 11 A2 10 VDD P L=1.8e-07 W=1.37e-06 $X=1965 $Y=2205 $D=16
M8 VDD A1 11 VDD P L=1.8e-07 W=1.37e-06 $X=2595 $Y=2205 $D=16
M9 Z 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3315 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INR4D2BWP7T A1 VDD B1 B2 ZN B3 VSS
** N=11 EP=7 IP=0 FDC=26
M0 8 A1 VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 ZN 8 VSS VSS N L=1.8e-07 W=1e-06 $X=2760 $Y=345 $D=0
M2 VSS 8 ZN VSS N L=1.8e-07 W=1e-06 $X=3480 $Y=345 $D=0
M3 ZN B1 VSS VSS N L=1.8e-07 W=1e-06 $X=5640 $Y=345 $D=0
M4 VSS B1 ZN VSS N L=1.8e-07 W=1e-06 $X=6360 $Y=345 $D=0
M5 ZN B2 VSS VSS N L=1.8e-07 W=1e-06 $X=9440 $Y=345 $D=0
M6 VSS B2 ZN VSS N L=1.8e-07 W=1e-06 $X=10160 $Y=345 $D=0
M7 ZN B3 VSS VSS N L=1.8e-07 W=1e-06 $X=12320 $Y=345 $D=0
M8 VSS B3 ZN VSS N L=1.8e-07 W=1e-06 $X=13040 $Y=345 $D=0
M9 8 A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M10 VDD 8 9 VDD P L=1.8e-07 W=1.37e-06 $X=2040 $Y=2205 $D=16
M11 9 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2760 $Y=2205 $D=16
M12 VDD 8 9 VDD P L=1.8e-07 W=1.37e-06 $X=3480 $Y=2205 $D=16
M13 9 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4200 $Y=2205 $D=16
M14 10 B1 9 VDD P L=1.8e-07 W=1.37e-06 $X=4920 $Y=2205 $D=16
M15 9 B1 10 VDD P L=1.8e-07 W=1.37e-06 $X=5640 $Y=2205 $D=16
M16 10 B1 9 VDD P L=1.8e-07 W=1.37e-06 $X=6360 $Y=2205 $D=16
M17 9 B1 10 VDD P L=1.8e-07 W=1.37e-06 $X=7080 $Y=2205 $D=16
M18 10 B2 11 VDD P L=1.8e-07 W=1.37e-06 $X=8720 $Y=2205 $D=16
M19 11 B2 10 VDD P L=1.8e-07 W=1.37e-06 $X=9440 $Y=2205 $D=16
M20 10 B2 11 VDD P L=1.8e-07 W=1.37e-06 $X=10160 $Y=2205 $D=16
M21 11 B2 10 VDD P L=1.8e-07 W=1.37e-06 $X=10880 $Y=2205 $D=16
M22 ZN B3 11 VDD P L=1.8e-07 W=1.37e-06 $X=11600 $Y=2205 $D=16
M23 11 B3 ZN VDD P L=1.8e-07 W=1.37e-06 $X=12320 $Y=2205 $D=16
M24 ZN B3 11 VDD P L=1.8e-07 W=1.37e-06 $X=13040 $Y=2205 $D=16
M25 11 B3 ZN VDD P L=1.8e-07 W=1.37e-06 $X=13760 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AO211D2BWP7T A1 A2 B C Z VSS VDD
** N=11 EP=7 IP=0 FDC=12
M0 10 A1 9 VSS N L=1.8e-07 W=1e-06 $X=660 $Y=345 $D=0
M1 VSS A2 10 VSS N L=1.8e-07 W=1e-06 $X=1140 $Y=345 $D=0
M2 9 B VSS VSS N L=1.8e-07 W=1e-06 $X=2020 $Y=345 $D=0
M3 VSS C 9 VSS N L=1.8e-07 W=1e-06 $X=2740 $Y=345 $D=0
M4 Z 9 VSS VSS N L=1.8e-07 W=1e-06 $X=3460 $Y=345 $D=0
M5 VSS 9 Z VSS N L=1.8e-07 W=1e-06 $X=4180 $Y=345 $D=0
M6 9 A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M7 8 A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=1380 $Y=2205 $D=16
M8 11 B 8 VDD P L=1.8e-07 W=1.37e-06 $X=2100 $Y=2205 $D=16
M9 VDD C 11 VDD P L=1.8e-07 W=1.37e-06 $X=2700 $Y=2205 $D=16
M10 Z 9 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3460 $Y=2205 $D=16
M11 VDD 9 Z VDD P L=1.8e-07 W=1.37e-06 $X=4180 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OAI211D0BWP7T C VSS B A1 VDD A2 ZN
** N=10 EP=7 IP=0 FDC=8
M0 8 C VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=680 $D=0
M1 9 B 8 VSS N L=1.8e-07 W=5e-07 $X=1115 $Y=680 $D=0
M2 ZN A1 9 VSS N L=1.8e-07 W=5e-07 $X=1820 $Y=680 $D=0
M3 9 A2 ZN VSS N L=1.8e-07 W=5e-07 $X=2560 $Y=680 $D=0
M4 ZN C VDD VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2830 $D=16
M5 VDD B ZN VDD P L=1.8e-07 W=6.85e-07 $X=1340 $Y=2830 $D=16
M6 10 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=2060 $Y=2830 $D=16
M7 ZN A2 10 VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2830 $D=16
.ENDS
***************************************
.SUBCKT CKND2D1BWP7T A2 VSS A1 ZN VDD
** N=6 EP=5 IP=0 FDC=4
M0 6 A2 VSS VSS N L=1.8e-07 W=6.85e-07 $X=660 $Y=345 $D=0
M1 ZN A1 6 VSS N L=1.8e-07 W=1e-06 $X=1385 $Y=345 $D=0
M2 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M3 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1385 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OAI211D2BWP7T C VSS B A2 ZN A1 VDD
** N=12 EP=7 IP=0 FDC=16
M0 9 B 8 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS C 9 VSS N L=1.8e-07 W=1e-06 $X=1120 $Y=345 $D=0
M2 10 C VSS VSS N L=1.8e-07 W=1e-06 $X=1950 $Y=345 $D=0
M3 8 B 10 VSS N L=1.8e-07 W=1e-06 $X=2480 $Y=345 $D=0
M4 ZN A1 8 VSS N L=1.8e-07 W=1e-06 $X=3200 $Y=345 $D=0
M5 8 A2 ZN VSS N L=1.8e-07 W=1e-06 $X=3920 $Y=345 $D=0
M6 ZN A2 8 VSS N L=1.8e-07 W=1e-06 $X=4640 $Y=345 $D=0
M7 8 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=5360 $Y=345 $D=0
M8 ZN B VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M9 VDD C ZN VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M10 ZN C VDD VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M11 VDD B ZN VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M12 11 A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3560 $Y=2205 $D=16
M13 ZN A2 11 VDD P L=1.8e-07 W=1.37e-06 $X=4020 $Y=2205 $D=16
M14 12 A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4740 $Y=2205 $D=16
M15 VDD A1 12 VDD P L=1.8e-07 W=1.37e-06 $X=5320 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKND2D0BWP7T A2 VSS A1 ZN VDD
** N=6 EP=5 IP=0 FDC=4
M0 6 A2 VSS VSS N L=1.8e-07 W=4.2e-07 $X=660 $Y=575 $D=0
M1 ZN A1 6 VSS N L=1.8e-07 W=4.8e-07 $X=1315 $Y=575 $D=0
M2 ZN A2 VDD VDD P L=1.8e-07 W=8e-07 $X=660 $Y=2765 $D=16
M3 VDD A1 ZN VDD P L=1.8e-07 W=8e-07 $X=1385 $Y=2765 $D=16
.ENDS
***************************************
.SUBCKT CKND2D3BWP7T A2 VSS ZN A1 VDD
** N=6 EP=5 IP=0 FDC=12
M0 6 A2 VSS VSS N L=1.8e-07 W=6e-07 $X=620 $Y=450 $D=0
M1 VSS A2 6 VSS N L=1.8e-07 W=6e-07 $X=1340 $Y=450 $D=0
M2 6 A2 VSS VSS N L=1.8e-07 W=6e-07 $X=2060 $Y=450 $D=0
M3 ZN A1 6 VSS N L=1.8e-07 W=8e-07 $X=2780 $Y=450 $D=0
M4 6 A1 ZN VSS N L=1.8e-07 W=8e-07 $X=3520 $Y=450 $D=0
M5 ZN A1 6 VSS N L=1.8e-07 W=8e-07 $X=4240 $Y=450 $D=0
M6 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M7 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M8 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M9 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M10 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3505 $Y=2205 $D=16
M11 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4225 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AO211D0BWP7T A1 A2 B C VSS VDD Z
** N=11 EP=7 IP=0 FDC=10
M0 9 A1 8 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=845 $D=0
M1 VSS A2 9 VSS N L=1.8e-07 W=5e-07 $X=1050 $Y=845 $D=0
M2 8 B VSS VSS N L=1.8e-07 W=5e-07 $X=1780 $Y=880 $D=0
M3 VSS C 8 VSS N L=1.8e-07 W=5e-07 $X=2500 $Y=880 $D=0
M4 Z 8 VSS VSS N L=1.8e-07 W=5e-07 $X=3120 $Y=580 $D=0
M5 8 A1 10 VDD P L=1.8e-07 W=6.85e-07 $X=570 $Y=2395 $D=16
M6 10 A2 8 VDD P L=1.8e-07 W=6.85e-07 $X=1290 $Y=2395 $D=16
M7 11 B 10 VDD P L=1.8e-07 W=6.85e-07 $X=1970 $Y=2790 $D=16
M8 VDD C 11 VDD P L=1.8e-07 W=6.85e-07 $X=2400 $Y=2790 $D=16
M9 Z 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=3120 $Y=2790 $D=16
.ENDS
***************************************
.SUBCKT AOI211D2BWP7T C VDD B ZN A1 A2 VSS
** N=12 EP=7 IP=0 FDC=16
M0 ZN B VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS C ZN VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 ZN C VSS VSS N L=1.8e-07 W=1e-06 $X=2060 $Y=345 $D=0
M3 VSS B ZN VSS N L=1.8e-07 W=1e-06 $X=2780 $Y=345 $D=0
M4 9 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=3580 $Y=345 $D=0
M5 ZN A1 9 VSS N L=1.8e-07 W=1e-06 $X=4020 $Y=345 $D=0
M6 10 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=4740 $Y=345 $D=0
M7 VSS A2 10 VSS N L=1.8e-07 W=1e-06 $X=5320 $Y=345 $D=0
M8 11 B 8 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M9 VDD C 11 VDD P L=1.8e-07 W=1.37e-06 $X=1120 $Y=2205 $D=16
M10 12 C VDD VDD P L=1.8e-07 W=1.37e-06 $X=1920 $Y=2205 $D=16
M11 8 B 12 VDD P L=1.8e-07 W=1.37e-06 $X=2480 $Y=2205 $D=16
M12 ZN A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=3200 $Y=2205 $D=16
M13 8 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3920 $Y=2205 $D=16
M14 ZN A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=4640 $Y=2205 $D=16
M15 8 A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=5360 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR2D3BWP7T A2 VDD ZN A1 VSS
** N=6 EP=5 IP=0 FDC=12
M0 ZN A2 VSS VSS N L=1.8e-07 W=1e-06 $X=640 $Y=345 $D=0
M1 VSS A2 ZN VSS N L=1.8e-07 W=1e-06 $X=1360 $Y=345 $D=0
M2 ZN A2 VSS VSS N L=1.8e-07 W=1e-06 $X=2080 $Y=345 $D=0
M3 VSS A1 ZN VSS N L=1.8e-07 W=1e-06 $X=2800 $Y=345 $D=0
M4 ZN A1 VSS VSS N L=1.8e-07 W=1e-06 $X=3520 $Y=345 $D=0
M5 VSS A1 ZN VSS N L=1.8e-07 W=1e-06 $X=4240 $Y=345 $D=0
M6 6 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=640 $Y=2205 $D=16
M7 VDD A2 6 VDD P L=1.8e-07 W=1.37e-06 $X=1360 $Y=2205 $D=16
M8 6 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2080 $Y=2205 $D=16
M9 ZN A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=2800 $Y=2205 $D=16
M10 6 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3520 $Y=2205 $D=16
M11 ZN A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=4240 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT MOAI22D0BWP7T B1 B2 VSS VDD A1 ZN A2
** N=11 EP=7 IP=0 FDC=10
M0 9 B1 8 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=610 $D=0
M1 VSS B2 9 VSS N L=1.8e-07 W=5e-07 $X=1050 $Y=610 $D=0
M2 10 8 VSS VSS N L=1.8e-07 W=5e-07 $X=1850 $Y=610 $D=0
M3 ZN A1 10 VSS N L=1.8e-07 W=5e-07 $X=2560 $Y=845 $D=0
M4 10 A2 ZN VSS N L=1.8e-07 W=5e-07 $X=3280 $Y=845 $D=0
M5 8 B1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=460 $Y=2390 $D=16
M6 VDD B2 8 VDD P L=1.8e-07 W=6.85e-07 $X=1180 $Y=2390 $D=16
M7 ZN 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1980 $Y=2390 $D=16
M8 11 A1 ZN VDD P L=1.8e-07 W=6.85e-07 $X=2700 $Y=2390 $D=16
M9 VDD A2 11 VDD P L=1.8e-07 W=6.85e-07 $X=3280 $Y=2390 $D=16
.ENDS
***************************************
.SUBCKT AN2D1BWP7T A1 A2 VSS VDD Z
** N=7 EP=5 IP=0 FDC=6
M0 7 A1 6 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=345 $D=0
M1 VSS A2 7 VSS N L=1.8e-07 W=5e-07 $X=1205 $Y=345 $D=0
M2 Z 6 VSS VSS N L=1.8e-07 W=1e-06 $X=2000 $Y=345 $D=0
M3 6 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=520 $Y=2205 $D=16
M4 VDD A2 6 VDD P L=1.8e-07 W=6.85e-07 $X=1240 $Y=2205 $D=16
M5 Z 6 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2000 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ND2D2BWP7T A1 ZN A2 VSS VDD
** N=7 EP=5 IP=0 FDC=8
M0 6 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=700 $Y=345 $D=0
M1 ZN A1 6 VSS N L=1.8e-07 W=1e-06 $X=1420 $Y=345 $D=0
M2 7 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=2260 $Y=345 $D=0
M3 VSS A2 7 VSS N L=1.8e-07 W=1e-06 $X=2980 $Y=345 $D=0
M4 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=700 $Y=2205 $D=16
M5 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1420 $Y=2205 $D=16
M6 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2260 $Y=2205 $D=16
M7 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2980 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AOI221D1BWP7T C VDD B1 B2 A2 VSS A1 ZN
** N=12 EP=8 IP=0 FDC=10
M0 ZN C VSS VSS N L=1.8e-07 W=1e-06 $X=625 $Y=345 $D=0
M1 11 B1 ZN VSS N L=1.8e-07 W=1e-06 $X=1345 $Y=345 $D=0
M2 VSS B2 11 VSS N L=1.8e-07 W=1e-06 $X=2065 $Y=345 $D=0
M3 12 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=3520 $Y=345 $D=0
M4 ZN A1 12 VSS N L=1.8e-07 W=1e-06 $X=4240 $Y=345 $D=0
M5 9 C VDD VDD P L=1.8e-07 W=1.37e-06 $X=625 $Y=2205 $D=16
M6 10 B1 9 VDD P L=1.8e-07 W=1.37e-06 $X=1345 $Y=2205 $D=16
M7 9 B2 10 VDD P L=1.8e-07 W=1.37e-06 $X=2065 $Y=2205 $D=16
M8 ZN A2 10 VDD P L=1.8e-07 W=1.37e-06 $X=3520 $Y=2205 $D=16
M9 10 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4240 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR3D0BWP7T A3 VSS VDD A2 A1 ZN
** N=8 EP=6 IP=0 FDC=6
M0 ZN A3 VSS VSS N L=1.8e-07 W=5e-07 $X=625 $Y=770 $D=0
M1 VSS A2 ZN VSS N L=1.8e-07 W=5e-07 $X=1345 $Y=770 $D=0
M2 ZN A1 VSS VSS N L=1.8e-07 W=5e-07 $X=2000 $Y=770 $D=0
M3 7 A3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=625 $Y=2205 $D=16
M4 8 A2 7 VDD P L=1.8e-07 W=1.37e-06 $X=1225 $Y=2205 $D=16
M5 ZN A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=1825 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AOI21D1BWP7T A1 A2 VSS B ZN VDD
** N=8 EP=6 IP=0 FDC=6
M0 8 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=760 $Y=345 $D=0
M1 VSS A2 8 VSS N L=1.8e-07 W=1e-06 $X=1480 $Y=345 $D=0
M2 ZN B VSS VSS N L=1.8e-07 W=1e-06 $X=2200 $Y=345 $D=0
M3 ZN A1 7 VDD P L=1.8e-07 W=1.37e-06 $X=760 $Y=2205 $D=16
M4 7 A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1480 $Y=2205 $D=16
M5 VDD B 7 VDD P L=1.8e-07 W=1.37e-06 $X=2200 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ND3D2BWP7T A1 A2 ZN A3 VDD VSS
** N=10 EP=6 IP=0 FDC=12
M0 7 A3 VSS VSS N L=1.8e-07 W=1e-06 $X=700 $Y=345 $D=0
M1 8 A2 7 VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 ZN A1 8 VSS N L=1.8e-07 W=1e-06 $X=1980 $Y=345 $D=0
M3 9 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=2780 $Y=345 $D=0
M4 10 A2 9 VSS N L=1.8e-07 W=1e-06 $X=3500 $Y=345 $D=0
M5 VSS A3 10 VSS N L=1.8e-07 W=1e-06 $X=4220 $Y=345 $D=0
M6 ZN A3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M7 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M8 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M9 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M10 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3500 $Y=2205 $D=16
M11 VDD A3 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4220 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR2D0BWP7T A2 VDD A1 ZN VSS
** N=6 EP=5 IP=0 FDC=4
M0 ZN A2 VSS VSS N L=1.8e-07 W=5e-07 $X=660 $Y=500 $D=0
M1 VSS A1 ZN VSS N L=1.8e-07 W=5e-07 $X=1380 $Y=500 $D=0
M2 6 A2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=660 $Y=2735 $D=16
M3 ZN A1 6 VDD P L=1.8e-07 W=6.85e-07 $X=1260 $Y=2735 $D=16
.ENDS
***************************************
.SUBCKT ND4D2BWP7T A1 A2 A3 A4 ZN VSS VDD
** N=10 EP=7 IP=0 FDC=16
M0 ZN A1 8 VSS N L=1.8e-07 W=1e-06 $X=665 $Y=345 $D=0
M1 8 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=1385 $Y=345 $D=0
M2 9 A2 8 VSS N L=1.8e-07 W=1e-06 $X=2105 $Y=345 $D=0
M3 8 A2 9 VSS N L=1.8e-07 W=1e-06 $X=2825 $Y=345 $D=0
M4 9 A3 10 VSS N L=1.8e-07 W=1e-06 $X=4305 $Y=345 $D=0
M5 10 A3 9 VSS N L=1.8e-07 W=1e-06 $X=5025 $Y=345 $D=0
M6 VSS A4 10 VSS N L=1.8e-07 W=1e-06 $X=5745 $Y=345 $D=0
M7 10 A4 VSS VSS N L=1.8e-07 W=1e-06 $X=6465 $Y=345 $D=0
M8 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=665 $Y=2205 $D=16
M9 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1385 $Y=2205 $D=16
M10 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2345 $Y=2205 $D=16
M11 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3065 $Y=2205 $D=16
M12 ZN A3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3985 $Y=2205 $D=16
M13 VDD A3 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4705 $Y=2205 $D=16
M14 ZN A4 VDD VDD P L=1.8e-07 W=1.37e-06 $X=5645 $Y=2205 $D=16
M15 VDD A4 ZN VDD P L=1.8e-07 W=1.37e-06 $X=6365 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OAI31D2BWP7T B VSS ZN A3 A1 A2 VDD
** N=12 EP=7 IP=0 FDC=16
M0 VSS B 8 VSS N L=1.8e-07 W=9.3e-07 $X=620 $Y=345 $D=0
M1 8 B VSS VSS N L=1.8e-07 W=9.3e-07 $X=1420 $Y=345 $D=0
M2 ZN A1 8 VSS N L=1.8e-07 W=9.3e-07 $X=2140 $Y=345 $D=0
M3 8 A1 ZN VSS N L=1.8e-07 W=9.3e-07 $X=2860 $Y=345 $D=0
M4 ZN A3 8 VSS N L=1.8e-07 W=9.3e-07 $X=3580 $Y=345 $D=0
M5 8 A3 ZN VSS N L=1.8e-07 W=9.3e-07 $X=4300 $Y=345 $D=0
M6 ZN A2 8 VSS N L=1.8e-07 W=9.3e-07 $X=5020 $Y=345 $D=0
M7 8 A2 ZN VSS N L=1.8e-07 W=9.3e-07 $X=5740 $Y=345 $D=0
M8 ZN B VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M9 VDD B ZN VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M10 9 A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2140 $Y=2205 $D=16
M11 10 A2 9 VDD P L=1.8e-07 W=1.25e-06 $X=2860 $Y=2325 $D=16
M12 ZN A3 10 VDD P L=1.8e-07 W=1.305e-06 $X=3580 $Y=2270 $D=16
M13 11 A3 ZN VDD P L=1.8e-07 W=1.305e-06 $X=4300 $Y=2270 $D=16
M14 12 A2 11 VDD P L=1.8e-07 W=1.25e-06 $X=5020 $Y=2325 $D=16
M15 VDD A1 12 VDD P L=1.8e-07 W=1.25e-06 $X=5740 $Y=2325 $D=16
.ENDS
***************************************
.SUBCKT ND3D1BWP7T A3 VSS A2 A1 VDD ZN
** N=8 EP=6 IP=0 FDC=6
M0 7 A3 VSS VSS N L=1.8e-07 W=1e-06 $X=750 $Y=345 $D=0
M1 8 A2 7 VSS N L=1.8e-07 W=1e-06 $X=1350 $Y=345 $D=0
M2 ZN A1 8 VSS N L=1.8e-07 W=1e-06 $X=1950 $Y=345 $D=0
M3 ZN A3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=750 $Y=2205 $D=16
M4 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1470 $Y=2205 $D=16
M5 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2190 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AOI211D1BWP7T C VDD B A2 VSS ZN A1
** N=10 EP=7 IP=0 FDC=8
M0 ZN C VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS B ZN VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 9 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=2060 $Y=345 $D=0
M3 ZN A1 9 VSS N L=1.8e-07 W=1e-06 $X=2560 $Y=345 $D=0
M4 10 C VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M5 8 B 10 VDD P L=1.8e-07 W=1.37e-06 $X=1120 $Y=2205 $D=16
M6 ZN A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=1840 $Y=2205 $D=16
M7 8 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2560 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IND4D2BWP7T A1 VSS B1 B2 ZN B3 VDD
** N=11 EP=7 IP=0 FDC=18
M0 VSS A1 8 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS 8 9 VSS N L=1.8e-07 W=1e-06 $X=1920 $Y=345 $D=0
M2 9 8 VSS VSS N L=1.8e-07 W=1e-06 $X=2640 $Y=345 $D=0
M3 10 B1 9 VSS N L=1.8e-07 W=1e-06 $X=3360 $Y=345 $D=0
M4 9 B1 10 VSS N L=1.8e-07 W=1e-06 $X=4080 $Y=345 $D=0
M5 10 B2 11 VSS N L=1.8e-07 W=1e-06 $X=5440 $Y=345 $D=0
M6 11 B2 10 VSS N L=1.8e-07 W=1e-06 $X=6160 $Y=345 $D=0
M7 ZN B3 11 VSS N L=1.8e-07 W=1e-06 $X=6880 $Y=345 $D=0
M8 11 B3 ZN VSS N L=1.8e-07 W=1e-06 $X=7600 $Y=345 $D=0
M9 VDD A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M10 ZN 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1860 $Y=2205 $D=16
M11 VDD 8 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2580 $Y=2205 $D=16
M12 ZN B1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3300 $Y=2205 $D=16
M13 VDD B1 ZN VDD P L=1.8e-07 W=1.29e-06 $X=4020 $Y=2285 $D=16
M14 ZN B2 VDD VDD P L=1.8e-07 W=1.29e-06 $X=5440 $Y=2285 $D=16
M15 VDD B2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=6160 $Y=2205 $D=16
M16 ZN B3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=6880 $Y=2205 $D=16
M17 VDD B3 ZN VDD P L=1.8e-07 W=1.37e-06 $X=7600 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INR2D1BWP7T A1 VDD ZN B1 VSS
** N=7 EP=5 IP=0 FDC=6
M0 VSS A1 6 VSS N L=1.8e-07 W=5e-07 $X=640 $Y=845 $D=0
M1 ZN 6 VSS VSS N L=1.8e-07 W=1e-06 $X=1280 $Y=345 $D=0
M2 VSS B1 ZN VSS N L=1.8e-07 W=1e-06 $X=2000 $Y=345 $D=0
M3 VDD A1 6 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2890 $D=16
M4 7 6 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1420 $Y=2205 $D=16
M5 ZN B1 7 VDD P L=1.8e-07 W=1.37e-06 $X=2000 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456
** N=1182 EP=456 IP=6778 FDC=10593
M0 28 5 1 1 N L=1.8e-07 W=1e-06 $X=38790 $Y=473375 $D=0
M1 1 5 28 1 N L=1.8e-07 W=1e-06 $X=39510 $Y=473375 $D=0
M2 28 5 1 1 N L=1.8e-07 W=1e-06 $X=40270 $Y=473375 $D=0
M3 1 5 28 1 N L=1.8e-07 W=1e-06 $X=40990 $Y=473375 $D=0
M4 28 5 1 1 N L=1.8e-07 W=1e-06 $X=41770 $Y=473375 $D=0
M5 1 5 28 1 N L=1.8e-07 W=1e-06 $X=42490 $Y=473375 $D=0
M6 28 5 1 1 N L=1.8e-07 W=1e-06 $X=43270 $Y=473375 $D=0
M7 1 5 28 1 N L=1.8e-07 W=1e-06 $X=43990 $Y=473375 $D=0
M8 28 5 1 1 N L=1.8e-07 W=1e-06 $X=44770 $Y=473375 $D=0
M9 1 5 28 1 N L=1.8e-07 W=1e-06 $X=45490 $Y=473375 $D=0
M10 1170 650 1 1 N L=1.8e-07 W=5e-07 $X=107460 $Y=459500 $D=0
M11 1171 689 1170 1 N L=1.8e-07 W=5e-07 $X=108130 $Y=459500 $D=0
M12 704 79 1171 1 N L=1.8e-07 W=5e-07 $X=108800 $Y=459500 $D=0
M13 1 687 704 1 N L=1.8e-07 W=5e-07 $X=109520 $Y=459500 $D=0
M14 713 704 1 1 N L=1.8e-07 W=5e-07 $X=110470 $Y=459500 $D=0
M15 464 708 1 1 N L=1.8e-07 W=1e-06 $X=133785 $Y=426335 $D=0
M16 1 708 464 1 N L=1.8e-07 W=1e-06 $X=134505 $Y=426335 $D=0
M17 464 708 1 1 N L=1.8e-07 W=1e-06 $X=135225 $Y=426335 $D=0
M18 1 708 464 1 N L=1.8e-07 W=1e-06 $X=135945 $Y=426335 $D=0
M19 464 708 1 1 N L=1.8e-07 W=1e-06 $X=136665 $Y=426335 $D=0
M20 1 708 464 1 N L=1.8e-07 W=1e-06 $X=137385 $Y=426335 $D=0
M21 464 708 1 1 N L=1.8e-07 W=1e-06 $X=138105 $Y=426335 $D=0
M22 1 708 464 1 N L=1.8e-07 W=1e-06 $X=138825 $Y=426335 $D=0
M23 464 742 1 1 N L=1.8e-07 W=1e-06 $X=139545 $Y=426335 $D=0
M24 1 742 464 1 N L=1.8e-07 W=1e-06 $X=140265 $Y=426335 $D=0
M25 464 742 1 1 N L=1.8e-07 W=1e-06 $X=140985 $Y=426335 $D=0
M26 1 742 464 1 N L=1.8e-07 W=1e-06 $X=141705 $Y=426335 $D=0
M27 464 742 1 1 N L=1.8e-07 W=1e-06 $X=142425 $Y=426335 $D=0
M28 1 742 464 1 N L=1.8e-07 W=1e-06 $X=143145 $Y=426335 $D=0
M29 464 742 1 1 N L=1.8e-07 W=1e-06 $X=143865 $Y=426335 $D=0
M30 1 742 464 1 N L=1.8e-07 W=1e-06 $X=144585 $Y=426335 $D=0
M31 841 144 1 1 N L=1.8e-07 W=1e-06 $X=168500 $Y=473375 $D=0
M32 166 810 1 1 N L=1.8e-07 W=1e-06 $X=170460 $Y=473375 $D=0
M33 1 810 166 1 N L=1.8e-07 W=1e-06 $X=171200 $Y=473375 $D=0
M34 166 150 1 1 N L=1.8e-07 W=1e-06 $X=173360 $Y=473375 $D=0
M35 1 150 166 1 N L=1.8e-07 W=1e-06 $X=174080 $Y=473375 $D=0
M36 166 841 1 1 N L=1.8e-07 W=1e-06 $X=177135 $Y=473375 $D=0
M37 1 841 166 1 N L=1.8e-07 W=1e-06 $X=177855 $Y=473375 $D=0
M38 166 864 1 1 N L=1.8e-07 W=1e-06 $X=180435 $Y=473375 $D=0
M39 1 864 166 1 N L=1.8e-07 W=1e-06 $X=181155 $Y=473375 $D=0
M40 1 862 864 1 N L=1.8e-07 W=1e-06 $X=182715 $Y=473375 $D=0
M41 1172 893 1 1 N L=1.8e-07 W=1e-06 $X=195400 $Y=442015 $D=0
M42 1173 828 1172 1 N L=1.8e-07 W=1e-06 $X=196020 $Y=442015 $D=0
M43 912 911 1173 1 N L=1.8e-07 W=1e-06 $X=196640 $Y=442015 $D=0
M44 1 880 912 1 N L=1.8e-07 W=1e-06 $X=197475 $Y=442015 $D=0
M45 916 912 1 1 N L=1.8e-07 W=1e-06 $X=198385 $Y=442015 $D=0
M46 1 882 931 1 N L=1.8e-07 W=4.2e-07 $X=209350 $Y=434665 $D=0
M47 946 881 1 1 N L=1.8e-07 W=5e-07 $X=210075 $Y=434585 $D=0
M48 1 204 946 1 N L=1.8e-07 W=5e-07 $X=210795 $Y=434585 $D=0
M49 946 931 1 1 N L=1.8e-07 W=5e-07 $X=211520 $Y=434585 $D=0
M50 1 941 946 1 N L=1.8e-07 W=5e-07 $X=212240 $Y=434585 $D=0
M51 941 890 1 1 N L=1.8e-07 W=4.2e-07 $X=212960 $Y=434665 $D=0
M52 1 1000 1005 1 N L=1.8e-07 W=5e-07 $X=251900 $Y=465780 $D=0
M53 1174 1008 1 1 N L=1.8e-07 W=5e-07 $X=252660 $Y=465605 $D=0
M54 1010 1000 1174 1 N L=1.8e-07 W=5e-07 $X=253290 $Y=465605 $D=0
M55 1008 1005 1010 1 N L=1.8e-07 W=5e-07 $X=254010 $Y=465605 $D=0
M56 1 239 1008 1 N L=1.8e-07 W=5e-07 $X=254790 $Y=465795 $D=0
M57 1 1010 1013 1 N L=1.8e-07 W=5e-07 $X=256210 $Y=465535 $D=0
M58 1175 1022 1 1 N L=1.8e-07 W=5e-07 $X=256930 $Y=465535 $D=0
M59 1014 1013 1175 1 N L=1.8e-07 W=5e-07 $X=257410 $Y=465535 $D=0
M60 1022 1010 1014 1 N L=1.8e-07 W=5e-07 $X=258170 $Y=465940 $D=0
M61 1 1014 1015 1 N L=1.8e-07 W=5e-07 $X=259600 $Y=465750 $D=0
M62 1025 1019 1 1 N L=1.8e-07 W=5e-07 $X=260400 $Y=465750 $D=0
M63 1022 1027 1025 1 N L=1.8e-07 W=5e-07 $X=261165 $Y=465605 $D=0
M64 1176 218 1022 1 N L=1.8e-07 W=5e-07 $X=261885 $Y=465605 $D=0
M65 1 1025 1176 1 N L=1.8e-07 W=5e-07 $X=262600 $Y=465605 $D=0
M66 1027 218 1 1 N L=1.8e-07 W=5e-07 $X=263360 $Y=465785 $D=0
M67 1 1058 1087 1 N L=1.8e-07 W=1e-06 $X=337585 $Y=467225 $D=0
M68 315 1087 1 1 N L=1.8e-07 W=1e-06 $X=338305 $Y=467225 $D=0
M69 28 5 2 2 P L=1.8e-07 W=1.37e-06 $X=38790 $Y=471145 $D=16
M70 2 5 28 2 P L=1.8e-07 W=1.37e-06 $X=39510 $Y=471145 $D=16
M71 28 5 2 2 P L=1.8e-07 W=1.37e-06 $X=40270 $Y=471145 $D=16
M72 2 5 28 2 P L=1.8e-07 W=1.37e-06 $X=40990 $Y=471145 $D=16
M73 28 5 2 2 P L=1.8e-07 W=1.37e-06 $X=41770 $Y=471145 $D=16
M74 2 5 28 2 P L=1.8e-07 W=1.37e-06 $X=42490 $Y=471145 $D=16
M75 28 5 2 2 P L=1.8e-07 W=1.37e-06 $X=43270 $Y=471145 $D=16
M76 2 5 28 2 P L=1.8e-07 W=1.37e-06 $X=43990 $Y=471145 $D=16
M77 28 5 2 2 P L=1.8e-07 W=1.37e-06 $X=44770 $Y=471145 $D=16
M78 2 5 28 2 P L=1.8e-07 W=1.37e-06 $X=45490 $Y=471145 $D=16
M79 703 650 704 2 P L=1.8e-07 W=6.85e-07 $X=107460 $Y=461655 $D=16
M80 704 689 703 2 P L=1.8e-07 W=6.85e-07 $X=108180 $Y=461655 $D=16
M81 703 79 704 2 P L=1.8e-07 W=6.85e-07 $X=108965 $Y=461655 $D=16
M82 2 687 703 2 P L=1.8e-07 W=6.85e-07 $X=109710 $Y=461655 $D=16
M83 713 704 2 2 P L=1.8e-07 W=6.85e-07 $X=110470 $Y=461655 $D=16
M84 2 708 773 2 P L=1.8e-07 W=1.37e-06 $X=133785 $Y=424105 $D=16
M85 773 708 2 2 P L=1.8e-07 W=1.37e-06 $X=134505 $Y=424105 $D=16
M86 2 708 773 2 P L=1.8e-07 W=1.37e-06 $X=135225 $Y=424105 $D=16
M87 773 708 2 2 P L=1.8e-07 W=1.37e-06 $X=135945 $Y=424105 $D=16
M88 2 708 773 2 P L=1.8e-07 W=1.37e-06 $X=136665 $Y=424105 $D=16
M89 773 708 2 2 P L=1.8e-07 W=1.37e-06 $X=137385 $Y=424105 $D=16
M90 2 708 773 2 P L=1.8e-07 W=1.37e-06 $X=138105 $Y=424105 $D=16
M91 773 708 2 2 P L=1.8e-07 W=1.37e-06 $X=138825 $Y=424105 $D=16
M92 464 742 773 2 P L=1.8e-07 W=1.37e-06 $X=139545 $Y=424105 $D=16
M93 773 742 464 2 P L=1.8e-07 W=1.37e-06 $X=140265 $Y=424105 $D=16
M94 464 742 773 2 P L=1.8e-07 W=1.37e-06 $X=140985 $Y=424105 $D=16
M95 773 742 464 2 P L=1.8e-07 W=1.37e-06 $X=141705 $Y=424105 $D=16
M96 464 742 773 2 P L=1.8e-07 W=1.37e-06 $X=142425 $Y=424105 $D=16
M97 773 742 464 2 P L=1.8e-07 W=1.37e-06 $X=143145 $Y=424105 $D=16
M98 464 742 773 2 P L=1.8e-07 W=1.37e-06 $X=143865 $Y=424105 $D=16
M99 773 742 464 2 P L=1.8e-07 W=1.37e-06 $X=144585 $Y=424105 $D=16
M100 841 144 2 2 P L=1.8e-07 W=1.37e-06 $X=168500 $Y=471145 $D=16
M101 2 810 837 2 P L=1.8e-07 W=1.37e-06 $X=169760 $Y=471145 $D=16
M102 837 810 2 2 P L=1.8e-07 W=1.37e-06 $X=170480 $Y=471145 $D=16
M103 2 810 837 2 P L=1.8e-07 W=1.37e-06 $X=171200 $Y=471145 $D=16
M104 837 810 2 2 P L=1.8e-07 W=1.37e-06 $X=171920 $Y=471145 $D=16
M105 850 150 837 2 P L=1.8e-07 W=1.37e-06 $X=172640 $Y=471145 $D=16
M106 837 150 850 2 P L=1.8e-07 W=1.37e-06 $X=173360 $Y=471145 $D=16
M107 850 150 837 2 P L=1.8e-07 W=1.37e-06 $X=174080 $Y=471145 $D=16
M108 837 150 850 2 P L=1.8e-07 W=1.37e-06 $X=174800 $Y=471145 $D=16
M109 850 841 863 2 P L=1.8e-07 W=1.37e-06 $X=176415 $Y=471145 $D=16
M110 863 841 850 2 P L=1.8e-07 W=1.37e-06 $X=177135 $Y=471145 $D=16
M111 850 841 863 2 P L=1.8e-07 W=1.37e-06 $X=177855 $Y=471145 $D=16
M112 863 841 850 2 P L=1.8e-07 W=1.37e-06 $X=178575 $Y=471145 $D=16
M113 166 864 863 2 P L=1.8e-07 W=1.37e-06 $X=179295 $Y=471145 $D=16
M114 863 864 166 2 P L=1.8e-07 W=1.37e-06 $X=180015 $Y=471145 $D=16
M115 166 864 863 2 P L=1.8e-07 W=1.37e-06 $X=180735 $Y=471145 $D=16
M116 863 864 166 2 P L=1.8e-07 W=1.37e-06 $X=181455 $Y=471145 $D=16
M117 2 862 864 2 P L=1.8e-07 W=1.37e-06 $X=182715 $Y=471145 $D=16
M118 909 893 912 2 P L=1.8e-07 W=1.37e-06 $X=195400 $Y=439785 $D=16
M119 912 828 909 2 P L=1.8e-07 W=1.37e-06 $X=196120 $Y=439785 $D=16
M120 909 911 912 2 P L=1.8e-07 W=1.37e-06 $X=196880 $Y=439785 $D=16
M121 2 880 909 2 P L=1.8e-07 W=1.37e-06 $X=197625 $Y=439785 $D=16
M122 916 912 2 2 P L=1.8e-07 W=1.37e-06 $X=198385 $Y=439785 $D=16
M123 2 882 931 2 P L=1.8e-07 W=4.2e-07 $X=209345 $Y=432200 $D=16
M124 1177 881 2 2 P L=1.8e-07 W=1.37e-06 $X=210145 $Y=431945 $D=16
M125 1178 204 1177 2 P L=1.8e-07 W=1.37e-06 $X=210715 $Y=431945 $D=16
M126 1179 931 1178 2 P L=1.8e-07 W=1.37e-06 $X=211285 $Y=431945 $D=16
M127 946 941 1179 2 P L=1.8e-07 W=1.37e-06 $X=211855 $Y=431945 $D=16
M128 2 890 941 2 P L=1.8e-07 W=4.2e-07 $X=213115 $Y=432780 $D=16
M129 2 1000 1005 2 P L=1.8e-07 W=6.85e-07 $X=251900 $Y=463520 $D=16
M130 1180 1008 2 2 P L=1.8e-07 W=6.85e-07 $X=252660 $Y=463765 $D=16
M131 1010 1005 1180 2 P L=1.8e-07 W=6.85e-07 $X=253290 $Y=463765 $D=16
M132 1008 1000 1010 2 P L=1.8e-07 W=6.85e-07 $X=254030 $Y=463765 $D=16
M133 2 239 1008 2 P L=1.8e-07 W=6.85e-07 $X=254750 $Y=463765 $D=16
M134 2 1010 1013 2 P L=1.8e-07 W=6.85e-07 $X=256210 $Y=463790 $D=16
M135 1181 1022 2 2 P L=1.8e-07 W=6.85e-07 $X=256930 $Y=463790 $D=16
M136 1014 1010 1181 2 P L=1.8e-07 W=6.85e-07 $X=257420 $Y=463790 $D=16
M137 1022 1013 1014 2 P L=1.8e-07 W=6.85e-07 $X=258160 $Y=463790 $D=16
M138 2 1014 1015 2 P L=1.8e-07 W=6.85e-07 $X=259600 $Y=463990 $D=16
M139 1025 1019 2 2 P L=1.8e-07 W=6.85e-07 $X=260400 $Y=463990 $D=16
M140 1022 218 1025 2 P L=1.8e-07 W=6.85e-07 $X=261165 $Y=463810 $D=16
M141 1182 1027 1022 2 P L=1.8e-07 W=6.85e-07 $X=261885 $Y=463810 $D=16
M142 2 1025 1182 2 P L=1.8e-07 W=6.85e-07 $X=262570 $Y=463810 $D=16
M143 1027 218 2 2 P L=1.8e-07 W=6.85e-07 $X=263360 $Y=463475 $D=16
M144 2 1058 1087 2 P L=1.8e-07 W=1.37e-06 $X=337585 $Y=469085 $D=16
M145 315 1087 2 2 P L=1.8e-07 W=1.37e-06 $X=338305 $Y=469085 $D=16
X205 1 5 ANTENNABWP7T $T=22240 474720 0 180 $X=20830 $Y=470510
X206 1 455 ANTENNABWP7T $T=474160 419840 0 180 $X=472750 $Y=415630
X207 1 437 ANTENNABWP7T $T=473040 419840 0 0 $X=472750 $Y=419605
X208 1 405 ANTENNABWP7T $T=473040 427680 0 0 $X=472750 $Y=427445
X209 1 407 ANTENNABWP7T $T=474160 435520 0 180 $X=472750 $Y=431310
X210 1 362 ANTENNABWP7T $T=473040 435520 0 0 $X=472750 $Y=435285
X211 1 435 ANTENNABWP7T $T=474160 443360 0 180 $X=472750 $Y=439150
X212 1 442 ANTENNABWP7T $T=473040 443360 0 0 $X=472750 $Y=443125
X213 1 443 ANTENNABWP7T $T=474160 451200 0 180 $X=472750 $Y=446990
X214 1 454 ANTENNABWP7T $T=473040 451200 0 0 $X=472750 $Y=450965
X215 1 456 ANTENNABWP7T $T=474160 466880 0 180 $X=472750 $Y=462670
X216 1 426 ANTENNABWP7T $T=473040 466880 0 0 $X=472750 $Y=466645
X217 1 222 ANTENNABWP7T $T=474160 474720 0 180 $X=472750 $Y=470510
X218 1 324 350 ICV_1 $T=466320 466880 0 0 $X=466030 $Y=466645
X219 1 290 363 ICV_1 $T=468560 466880 0 0 $X=468270 $Y=466645
X220 1 449 423 ICV_1 $T=469680 459040 0 0 $X=469390 $Y=458805
X221 1 367 453 ICV_1 $T=470800 419840 0 0 $X=470510 $Y=419605
X222 1 270 353 ICV_1 $T=470800 427680 0 0 $X=470510 $Y=427445
X223 1 358 432 ICV_1 $T=470800 435520 0 0 $X=470510 $Y=435285
X224 1 409 335 ICV_1 $T=470800 443360 0 0 $X=470510 $Y=443125
X225 1 452 346 ICV_1 $T=470800 451200 0 0 $X=470510 $Y=450965
X226 1 361 311 ICV_1 $T=470800 466880 0 0 $X=470510 $Y=466645
X227 1 375 428 ICV_1 $T=471920 459040 0 0 $X=471630 $Y=458805
X228 1 421 393 ICV_2 $T=465200 474720 0 180 $X=463790 $Y=470510
X229 1 434 439 ICV_2 $T=467440 474720 0 180 $X=466030 $Y=470510
X230 1 394 284 ICV_2 $T=469680 466880 0 180 $X=468270 $Y=462670
X231 1 326 427 ICV_2 $T=469680 474720 0 180 $X=468270 $Y=470510
X232 1 419 279 ICV_2 $T=470800 427680 0 180 $X=469390 $Y=423470
X233 1 386 451 ICV_2 $T=470800 459040 0 180 $X=469390 $Y=454830
X234 1 406 400 ICV_2 $T=471920 419840 0 180 $X=470510 $Y=415630
X235 1 440 305 ICV_2 $T=471920 435520 0 180 $X=470510 $Y=431310
X236 1 313 441 ICV_2 $T=471920 443360 0 180 $X=470510 $Y=439150
X237 1 401 379 ICV_2 $T=471920 451200 0 180 $X=470510 $Y=446990
X238 1 415 273 ICV_2 $T=471920 466880 0 180 $X=470510 $Y=462670
X239 1 349 446 ICV_2 $T=471920 474720 0 180 $X=470510 $Y=470510
X240 1 373 371 ICV_2 $T=473040 427680 0 180 $X=471630 $Y=423470
X241 1 277 424 ICV_2 $T=473040 459040 0 180 $X=471630 $Y=454830
X333 539 1 2 546 CKBD1BWP7T $T=54720 427680 0 0 $X=54430 $Y=427445
X334 459 1 2 586 CKBD1BWP7T $T=67040 451200 1 0 $X=66750 $Y=446990
X335 750 1 2 761 CKBD1BWP7T $T=135920 459040 0 0 $X=135630 $Y=458805
X336 748 1 2 786 CKBD1BWP7T $T=148240 466880 0 0 $X=147950 $Y=466645
X337 952 1 2 972 CKBD1BWP7T $T=224400 466880 1 0 $X=224110 $Y=462670
X338 360 1 2 1121 CKBD1BWP7T $T=397440 419840 1 180 $X=394910 $Y=419605
X339 370 1 2 1123 CKBD1BWP7T $T=404720 435520 0 180 $X=402190 $Y=431310
X340 418 1 2 351 CKBD1BWP7T $T=461840 435520 1 180 $X=459310 $Y=435285
X341 447 1 2 323 CKBD1BWP7T $T=470800 419840 0 180 $X=468270 $Y=415630
X342 21 1 2 488 INVD0BWP7T $T=29520 419840 1 0 $X=29230 $Y=415630
X343 487 1 2 511 INVD0BWP7T $T=44640 466880 1 0 $X=44350 $Y=462670
X344 461 1 2 529 INVD0BWP7T $T=51360 435520 0 0 $X=51070 $Y=435285
X345 462 1 2 537 INVD0BWP7T $T=54720 466880 1 0 $X=54430 $Y=462670
X346 518 1 2 573 INVD0BWP7T $T=63680 427680 1 0 $X=63390 $Y=423470
X347 556 1 2 504 INVD0BWP7T $T=65360 443360 1 180 $X=63390 $Y=443125
X348 33 1 2 589 INVD0BWP7T $T=69280 443360 1 0 $X=68990 $Y=439150
X349 59 1 2 588 INVD0BWP7T $T=87200 419840 1 180 $X=85230 $Y=419605
X350 593 1 2 623 INVD0BWP7T $T=87760 427680 1 180 $X=85790 $Y=427445
X351 610 1 2 632 INVD0BWP7T $T=87200 443360 1 0 $X=86910 $Y=439150
X352 582 1 2 641 INVD0BWP7T $T=90000 435520 1 0 $X=89710 $Y=431310
X353 471 1 2 630 INVD0BWP7T $T=94480 474720 0 180 $X=92510 $Y=470510
X354 659 1 2 639 INVD0BWP7T $T=97280 435520 1 180 $X=95310 $Y=435285
X355 591 1 2 73 INVD0BWP7T $T=103440 419840 0 180 $X=101470 $Y=415630
X356 693 1 2 680 INVD0BWP7T $T=108480 427680 1 180 $X=106510 $Y=427445
X357 18 1 2 631 INVD0BWP7T $T=108480 435520 1 180 $X=106510 $Y=435285
X358 655 1 2 712 INVD0BWP7T $T=109600 466880 1 0 $X=109310 $Y=462670
X359 83 1 2 618 INVD0BWP7T $T=113520 427680 1 180 $X=111550 $Y=427445
X360 557 1 2 698 INVD0BWP7T $T=123600 451200 0 180 $X=121630 $Y=446990
X361 732 1 2 741 INVD0BWP7T $T=129200 435520 0 0 $X=128910 $Y=435285
X362 708 1 2 747 INVD0BWP7T $T=133680 427680 1 180 $X=131710 $Y=427445
X363 608 1 2 746 INVD0BWP7T $T=135920 451200 0 180 $X=133950 $Y=446990
X364 759 1 2 762 INVD0BWP7T $T=146000 451200 0 180 $X=144030 $Y=446990
X365 776 1 2 790 INVD0BWP7T $T=149360 435520 1 0 $X=149070 $Y=431310
X366 123 1 2 795 INVD0BWP7T $T=154400 419840 1 180 $X=152430 $Y=419605
X367 119 1 2 804 INVD0BWP7T $T=155520 451200 1 0 $X=155230 $Y=446990
X368 831 1 2 819 INVD0BWP7T $T=172880 443360 0 180 $X=170910 $Y=439150
X369 800 1 2 851 INVD0BWP7T $T=179040 451200 0 0 $X=178750 $Y=450965
X370 130 1 2 876 INVD0BWP7T $T=186320 443360 1 0 $X=186030 $Y=439150
X371 178 1 2 867 INVD0BWP7T $T=190240 443360 1 180 $X=188270 $Y=443125
X372 894 1 2 805 INVD0BWP7T $T=190800 466880 0 180 $X=188830 $Y=462670
X373 174 1 2 883 INVD0BWP7T $T=190240 459040 1 0 $X=189950 $Y=454830
X374 832 1 2 898 INVD0BWP7T $T=190800 466880 1 0 $X=190510 $Y=462670
X375 892 1 2 919 INVD0BWP7T $T=205920 427680 0 0 $X=205630 $Y=427445
X376 186 1 2 920 INVD0BWP7T $T=206480 419840 0 0 $X=206190 $Y=419605
X377 187 1 2 917 INVD0BWP7T $T=209280 427680 1 0 $X=208990 $Y=423470
X378 205 1 2 835 INVD0BWP7T $T=212080 443360 0 180 $X=210110 $Y=439150
X379 207 1 2 942 INVD0BWP7T $T=212080 419840 0 0 $X=211790 $Y=419605
X380 848 1 2 930 INVD0BWP7T $T=213760 443360 0 180 $X=211790 $Y=439150
X381 964 1 2 953 INVD0BWP7T $T=221600 459040 0 180 $X=219630 $Y=454830
X382 954 1 2 961 INVD0BWP7T $T=222720 459040 1 180 $X=220750 $Y=458805
X383 929 1 2 966 INVD0BWP7T $T=221600 443360 1 0 $X=221310 $Y=439150
X384 934 1 2 960 INVD0BWP7T $T=222720 435520 1 0 $X=222430 $Y=431310
X385 223 1 2 968 INVD0BWP7T $T=232240 443360 1 180 $X=230270 $Y=443125
X386 972 1 2 984 INVD0BWP7T $T=235040 451200 1 0 $X=234750 $Y=446990
X387 235 1 2 999 INVD0BWP7T $T=247920 466880 1 0 $X=247630 $Y=462670
X388 908 1 2 1024 INVD0BWP7T $T=263600 474720 0 180 $X=261630 $Y=470510
X389 973 1 2 1020 INVD0BWP7T $T=263600 435520 0 0 $X=263310 $Y=435285
X390 230 1 2 1033 INVD0BWP7T $T=269200 474720 1 0 $X=268910 $Y=470510
X391 338 1 2 334 INVD0BWP7T $T=362720 419840 0 180 $X=360750 $Y=415630
X392 369 1 2 1127 INVD0BWP7T $T=402480 443360 1 0 $X=402190 $Y=439150
X393 251 1 2 1165 INVD0BWP7T $T=457920 435520 0 0 $X=457630 $Y=435285
X394 430 1 2 1168 INVD0BWP7T $T=469680 459040 0 180 $X=467710 $Y=454830
X395 702 92 1 2 BUFFD1P5BWP7T $T=138720 474720 1 0 $X=138430 $Y=470510
X396 764 780 1 2 BUFFD1P5BWP7T $T=143760 466880 1 0 $X=143470 $Y=462670
X397 1034 246 1 2 BUFFD1P5BWP7T $T=272000 419840 0 180 $X=268910 $Y=415630
X398 1023 256 1 2 BUFFD1P5BWP7T $T=280400 451200 1 0 $X=280110 $Y=446990
X399 1107 337 1 2 BUFFD1P5BWP7T $T=365520 451200 1 180 $X=362430 $Y=450965
X400 1119 330 1 2 BUFFD1P5BWP7T $T=389040 474720 0 180 $X=385950 $Y=470510
X401 1134 376 1 2 BUFFD1P5BWP7T $T=409200 435520 1 180 $X=406110 $Y=435285
X402 1009 414 1 2 BUFFD1P5BWP7T $T=446720 435520 0 0 $X=446430 $Y=435285
X403 1163 410 1 2 BUFFD1P5BWP7T $T=450080 466880 0 180 $X=446990 $Y=462670
X404 443 436 1 2 BUFFD1P5BWP7T $T=468000 459040 0 180 $X=464910 $Y=454830
X405 448 327 1 2 BUFFD1P5BWP7T $T=470800 419840 1 180 $X=467710 $Y=419605
X406 1169 1 2 450 INVD3BWP7T $T=467440 427680 0 0 $X=467150 $Y=427445
X407 269 270 2 1 269 1055 270 MAOI22D0BWP7T $T=299440 419840 0 0 $X=299150 $Y=419605
X408 282 279 2 1 282 281 279 MAOI22D0BWP7T $T=312880 419840 0 180 $X=308670 $Y=415630
X409 298 305 2 1 298 1082 305 MAOI22D0BWP7T $T=337520 435520 0 180 $X=333310 $Y=431310
X410 306 309 2 1 309 1084 306 MAOI22D0BWP7T $T=338640 419840 0 180 $X=334430 $Y=415630
X411 312 313 2 1 312 1088 313 MAOI22D0BWP7T $T=336400 443360 1 0 $X=336110 $Y=439150
X412 323 335 2 1 323 1095 335 MAOI22D0BWP7T $T=364960 443360 1 180 $X=360750 $Y=443125
X413 340 343 2 1 343 1102 340 MAOI22D0BWP7T $T=379520 419840 1 180 $X=375310 $Y=419605
X414 354 353 2 1 354 1108 353 MAOI22D0BWP7T $T=392400 435520 1 180 $X=388190 $Y=435285
X415 1123 358 2 1 1123 1124 358 MAOI22D0BWP7T $T=399120 435520 1 180 $X=394910 $Y=435285
X416 351 379 2 1 351 1112 379 MAOI22D0BWP7T $T=419840 443360 0 180 $X=415630 $Y=439150
X417 408 405 2 1 408 1145 405 MAOI22D0BWP7T $T=450080 435520 0 180 $X=445870 $Y=431310
X418 411 406 2 1 411 1159 406 MAOI22D0BWP7T $T=450640 419840 0 180 $X=446430 $Y=415630
X419 413 409 2 1 413 1157 409 MAOI22D0BWP7T $T=451200 443360 0 180 $X=446990 $Y=439150
X420 420 419 2 1 420 1158 419 MAOI22D0BWP7T $T=464640 427680 1 180 $X=460430 $Y=427445
X421 431 437 2 1 431 1160 437 MAOI22D0BWP7T $T=469680 427680 0 180 $X=465470 $Y=423470
X422 444 440 2 1 444 1149 440 MAOI22D0BWP7T $T=470800 435520 0 180 $X=466590 $Y=431310
X423 438 441 2 1 438 1152 441 MAOI22D0BWP7T $T=470800 435520 1 180 $X=466590 $Y=435285
X504 218 220 220 218 967 1 2 MAOI22D2BWP7T $T=228880 419840 1 180 $X=222430 $Y=419605
X505 968 767 767 968 974 1 2 MAOI22D2BWP7T $T=223280 451200 0 0 $X=222990 $Y=450965
X506 92 225 225 92 985 1 2 MAOI22D2BWP7T $T=228880 419840 1 0 $X=228590 $Y=415630
X507 232 978 978 232 1053 1 2 MAOI22D2BWP7T $T=289920 427680 0 0 $X=289630 $Y=427445
X508 429 432 429 432 1051 1 2 MAOI22D2BWP7T $T=468000 419840 0 180 $X=461550 $Y=415630
X509 445 442 445 442 1081 1 2 MAOI22D2BWP7T $T=470800 443360 1 180 $X=464350 $Y=443125
X510 435 433 1137 433 1 435 2 IAO22D2BWP7T $T=470800 443360 0 180 $X=464350 $Y=439150
X511 478 1 2 479 BUFFD1BWP7T $T=30640 427680 1 180 $X=28110 $Y=427445
X512 479 1 2 489 BUFFD1BWP7T $T=28960 443360 0 0 $X=28670 $Y=443125
X513 535 1 2 540 BUFFD1BWP7T $T=52480 466880 1 0 $X=52190 $Y=462670
X514 533 1 2 543 BUFFD1BWP7T $T=53040 443360 1 0 $X=52750 $Y=439150
X515 743 1 2 749 BUFFD1BWP7T $T=130880 435520 0 0 $X=130590 $Y=435285
X516 769 1 2 778 BUFFD1BWP7T $T=144880 443360 1 0 $X=144590 $Y=439150
X517 799 1 2 775 BUFFD1BWP7T $T=155520 451200 0 180 $X=152990 $Y=446990
X518 944 1 2 935 BUFFD1BWP7T $T=215440 466880 1 180 $X=212910 $Y=466645
X519 932 1 2 952 BUFFD1BWP7T $T=214320 466880 1 0 $X=214030 $Y=462670
X520 971 1 2 973 BUFFD1BWP7T $T=224400 435520 1 0 $X=224110 $Y=431310
X521 274 1 2 1057 BUFFD1BWP7T $T=303360 419840 0 180 $X=300830 $Y=415630
X522 345 1 2 1105 BUFFD1BWP7T $T=379520 427680 0 180 $X=376990 $Y=423470
X523 352 1 2 1117 BUFFD1BWP7T $T=389040 427680 0 180 $X=386510 $Y=423470
X524 388 1 2 385 BUFFD1BWP7T $T=426560 419840 0 180 $X=424030 $Y=415630
X525 387 1 2 1140 BUFFD1BWP7T $T=424320 443360 1 0 $X=424030 $Y=439150
X526 395 1 2 1150 BUFFD1BWP7T $T=436640 427680 0 0 $X=436350 $Y=427445
X527 1167 1 2 1169 BUFFD1BWP7T $T=464640 435520 1 0 $X=464350 $Y=431310
X528 1 2 DCAP4BWP7T $T=26720 435520 0 0 $X=26430 $Y=435285
X529 1 2 DCAP4BWP7T $T=41280 435520 0 0 $X=40990 $Y=435285
X530 1 2 DCAP4BWP7T $T=51920 443360 0 0 $X=51630 $Y=443125
X531 1 2 DCAP4BWP7T $T=55280 419840 0 0 $X=54990 $Y=419605
X532 1 2 DCAP4BWP7T $T=65360 435520 0 0 $X=65070 $Y=435285
X533 1 2 DCAP4BWP7T $T=90000 459040 1 0 $X=89710 $Y=454830
X534 1 2 DCAP4BWP7T $T=126400 443360 1 0 $X=126110 $Y=439150
X535 1 2 DCAP4BWP7T $T=128640 419840 1 0 $X=128350 $Y=415630
X536 1 2 DCAP4BWP7T $T=148240 443360 0 0 $X=147950 $Y=443125
X537 1 2 DCAP4BWP7T $T=165600 474720 1 0 $X=165310 $Y=470510
X538 1 2 DCAP4BWP7T $T=171760 419840 1 0 $X=171470 $Y=415630
X539 1 2 DCAP4BWP7T $T=180160 459040 0 0 $X=179870 $Y=458805
X540 1 2 DCAP4BWP7T $T=212640 443360 0 0 $X=212350 $Y=443125
X541 1 2 DCAP4BWP7T $T=227200 427680 1 0 $X=226910 $Y=423470
X542 1 2 DCAP4BWP7T $T=251280 419840 1 0 $X=250990 $Y=415630
X543 1 2 DCAP4BWP7T $T=253520 443360 0 0 $X=253230 $Y=443125
X544 1 2 DCAP4BWP7T $T=266960 419840 1 0 $X=266670 $Y=415630
X545 1 2 DCAP4BWP7T $T=272000 435520 0 0 $X=271710 $Y=435285
X546 1 2 DCAP4BWP7T $T=287120 419840 1 0 $X=286830 $Y=415630
X547 1 2 DCAP4BWP7T $T=310080 435520 0 0 $X=309790 $Y=435285
X548 1 2 DCAP4BWP7T $T=317360 419840 1 0 $X=317070 $Y=415630
X549 1 2 DCAP4BWP7T $T=325760 419840 0 0 $X=325470 $Y=419605
X550 1 2 DCAP4BWP7T $T=342000 435520 1 0 $X=341710 $Y=431310
X551 1 2 DCAP4BWP7T $T=367760 427680 0 0 $X=367470 $Y=427445
X552 1 2 DCAP4BWP7T $T=371120 443360 0 0 $X=370830 $Y=443125
X553 1 2 DCAP4BWP7T $T=379520 427680 1 0 $X=379230 $Y=423470
X554 1 2 DCAP4BWP7T $T=399680 443360 0 0 $X=399390 $Y=443125
X555 1 2 DCAP4BWP7T $T=404160 435520 0 0 $X=403870 $Y=435285
X556 1 2 DCAP4BWP7T $T=417600 466880 1 0 $X=417310 $Y=462670
X557 1 2 DCAP4BWP7T $T=422080 435520 1 0 $X=421790 $Y=431310
X558 1 2 DCAP4BWP7T $T=431600 443360 0 0 $X=431310 $Y=443125
X559 1 2 DCAP4BWP7T $T=437200 443360 1 0 $X=436910 $Y=439150
X560 1 2 DCAP4BWP7T $T=439440 427680 1 0 $X=439150 $Y=423470
X561 1 2 DCAP4BWP7T $T=451760 459040 0 0 $X=451470 $Y=458805
X562 1 2 DCAP4BWP7T $T=451760 474720 1 0 $X=451470 $Y=470510
X563 1 2 DCAP4BWP7T $T=459600 419840 1 0 $X=459310 $Y=415630
X564 1 2 ICV_3 $T=23920 443360 1 0 $X=23630 $Y=439150
X565 1 2 ICV_3 $T=31200 419840 1 0 $X=30910 $Y=415630
X566 1 2 ICV_3 $T=31200 427680 1 0 $X=30910 $Y=423470
X567 1 2 ICV_3 $T=31200 435520 1 0 $X=30910 $Y=431310
X568 1 2 ICV_3 $T=31200 443360 0 0 $X=30910 $Y=443125
X569 1 2 ICV_3 $T=31200 459040 1 0 $X=30910 $Y=454830
X570 1 2 ICV_3 $T=31200 459040 0 0 $X=30910 $Y=458805
X571 1 2 ICV_3 $T=31200 466880 1 0 $X=30910 $Y=462670
X572 1 2 ICV_3 $T=31200 474720 1 0 $X=30910 $Y=470510
X573 1 2 ICV_3 $T=39600 466880 1 0 $X=39310 $Y=462670
X574 1 2 ICV_3 $T=44640 419840 0 0 $X=44350 $Y=419605
X575 1 2 ICV_3 $T=64240 451200 1 0 $X=63950 $Y=446990
X576 1 2 ICV_3 $T=73200 459040 1 0 $X=72910 $Y=454830
X577 1 2 ICV_3 $T=95600 466880 1 0 $X=95310 $Y=462670
X578 1 2 ICV_3 $T=115200 419840 1 0 $X=114910 $Y=415630
X579 1 2 ICV_3 $T=115200 419840 0 0 $X=114910 $Y=419605
X580 1 2 ICV_3 $T=115200 435520 0 0 $X=114910 $Y=435285
X581 1 2 ICV_3 $T=115200 451200 0 0 $X=114910 $Y=450965
X582 1 2 ICV_3 $T=115200 459040 0 0 $X=114910 $Y=458805
X583 1 2 ICV_3 $T=115200 466880 0 0 $X=114910 $Y=466645
X584 1 2 ICV_3 $T=115200 474720 1 0 $X=114910 $Y=470510
X585 1 2 ICV_3 $T=135920 474720 1 0 $X=135630 $Y=470510
X586 1 2 ICV_3 $T=142080 443360 1 0 $X=141790 $Y=439150
X587 1 2 ICV_3 $T=157200 419840 0 0 $X=156910 $Y=419605
X588 1 2 ICV_3 $T=157200 427680 1 0 $X=156910 $Y=423470
X589 1 2 ICV_3 $T=157200 451200 1 0 $X=156910 $Y=446990
X590 1 2 ICV_3 $T=157200 451200 0 0 $X=156910 $Y=450965
X591 1 2 ICV_3 $T=157200 459040 0 0 $X=156910 $Y=458805
X592 1 2 ICV_3 $T=157200 466880 1 0 $X=156910 $Y=462670
X593 1 2 ICV_3 $T=161120 466880 0 0 $X=160830 $Y=466645
X594 1 2 ICV_3 $T=180720 451200 1 0 $X=180430 $Y=446990
X595 1 2 ICV_3 $T=199200 435520 1 0 $X=198910 $Y=431310
X596 1 2 ICV_3 $T=199200 435520 0 0 $X=198910 $Y=435285
X597 1 2 ICV_3 $T=199200 459040 1 0 $X=198910 $Y=454830
X598 1 2 ICV_3 $T=199200 474720 1 0 $X=198910 $Y=470510
X599 1 2 ICV_3 $T=203120 427680 0 0 $X=202830 $Y=427445
X600 1 2 ICV_3 $T=208160 474720 1 0 $X=207870 $Y=470510
X601 1 2 ICV_3 $T=222720 459040 0 0 $X=222430 $Y=458805
X602 1 2 ICV_3 $T=226640 474720 1 0 $X=226350 $Y=470510
X603 1 2 ICV_3 $T=241200 451200 1 0 $X=240910 $Y=446990
X604 1 2 ICV_3 $T=245120 451200 0 0 $X=244830 $Y=450965
X605 1 2 ICV_3 $T=245120 474720 1 0 $X=244830 $Y=470510
X606 1 2 ICV_3 $T=251280 451200 0 0 $X=250990 $Y=450965
X607 1 2 ICV_3 $T=258560 427680 0 0 $X=258270 $Y=427445
X608 1 2 ICV_3 $T=264160 466880 1 0 $X=263870 $Y=462670
X609 1 2 ICV_3 $T=277600 451200 1 0 $X=277310 $Y=446990
X610 1 2 ICV_3 $T=283200 427680 1 0 $X=282910 $Y=423470
X611 1 2 ICV_3 $T=283200 451200 1 0 $X=282910 $Y=446990
X612 1 2 ICV_3 $T=283200 459040 1 0 $X=282910 $Y=454830
X613 1 2 ICV_3 $T=283200 466880 0 0 $X=282910 $Y=466645
X614 1 2 ICV_3 $T=294400 419840 1 0 $X=294110 $Y=415630
X615 1 2 ICV_3 $T=305600 451200 0 0 $X=305310 $Y=450965
X616 1 2 ICV_3 $T=310080 459040 0 0 $X=309790 $Y=458805
X617 1 2 ICV_3 $T=312880 459040 1 0 $X=312590 $Y=454830
X618 1 2 ICV_3 $T=325200 427680 1 0 $X=324910 $Y=423470
X619 1 2 ICV_3 $T=325200 459040 1 0 $X=324910 $Y=454830
X620 1 2 ICV_3 $T=325200 459040 0 0 $X=324910 $Y=458805
X621 1 2 ICV_3 $T=325200 466880 1 0 $X=324910 $Y=462670
X622 1 2 ICV_3 $T=325200 474720 1 0 $X=324910 $Y=470510
X623 1 2 ICV_3 $T=333600 443360 1 0 $X=333310 $Y=439150
X624 1 2 ICV_3 $T=340880 474720 1 0 $X=340590 $Y=470510
X625 1 2 ICV_3 $T=345920 451200 1 0 $X=345630 $Y=446990
X626 1 2 ICV_3 $T=367200 419840 1 0 $X=366910 $Y=415630
X627 1 2 ICV_3 $T=367200 419840 0 0 $X=366910 $Y=419605
X628 1 2 ICV_3 $T=367200 435520 1 0 $X=366910 $Y=431310
X629 1 2 ICV_3 $T=375600 466880 1 0 $X=375310 $Y=462670
X630 1 2 ICV_3 $T=375600 466880 0 0 $X=375310 $Y=466645
X631 1 2 ICV_3 $T=388480 419840 0 0 $X=388190 $Y=419605
X632 1 2 ICV_3 $T=389600 459040 1 0 $X=389310 $Y=454830
X633 1 2 ICV_3 $T=394640 443360 1 0 $X=394350 $Y=439150
X634 1 2 ICV_3 $T=409200 435520 0 0 $X=408910 $Y=435285
X635 1 2 ICV_3 $T=409200 459040 1 0 $X=408910 $Y=454830
X636 1 2 ICV_3 $T=409200 474720 1 0 $X=408910 $Y=470510
X637 1 2 ICV_3 $T=417600 435520 0 0 $X=417310 $Y=435285
X638 1 2 ICV_3 $T=432720 451200 0 0 $X=432430 $Y=450965
X639 1 2 ICV_3 $T=444480 466880 1 0 $X=444190 $Y=462670
X640 1 2 ICV_3 $T=451200 451200 1 0 $X=450910 $Y=446990
X641 1 2 ICV_3 $T=451200 466880 0 0 $X=450910 $Y=466645
X642 1 2 ICV_3 $T=455120 443360 1 0 $X=454830 $Y=439150
X643 1 2 ICV_3 $T=464640 427680 0 0 $X=464350 $Y=427445
X644 1 2 DCAP8BWP7T $T=35120 419840 0 0 $X=34830 $Y=419605
X645 1 2 DCAP8BWP7T $T=56960 419840 1 0 $X=56670 $Y=415630
X646 1 2 DCAP8BWP7T $T=70960 419840 1 0 $X=70670 $Y=415630
X647 1 2 DCAP8BWP7T $T=77120 466880 0 0 $X=76830 $Y=466645
X648 1 2 DCAP8BWP7T $T=112960 435520 1 0 $X=112670 $Y=431310
X649 1 2 DCAP8BWP7T $T=113520 427680 0 0 $X=113230 $Y=427445
X650 1 2 DCAP8BWP7T $T=113520 459040 1 0 $X=113230 $Y=454830
X651 1 2 DCAP8BWP7T $T=126960 427680 1 0 $X=126670 $Y=423470
X652 1 2 DCAP8BWP7T $T=137040 443360 0 0 $X=136750 $Y=443125
X653 1 2 DCAP8BWP7T $T=137040 451200 0 0 $X=136750 $Y=450965
X654 1 2 DCAP8BWP7T $T=147680 419840 0 0 $X=147390 $Y=419605
X655 1 2 DCAP8BWP7T $T=155520 443360 0 0 $X=155230 $Y=443125
X656 1 2 DCAP8BWP7T $T=168400 451200 1 0 $X=168110 $Y=446990
X657 1 2 DCAP8BWP7T $T=195840 466880 0 0 $X=195550 $Y=466645
X658 1 2 DCAP8BWP7T $T=216560 466880 1 0 $X=216270 $Y=462670
X659 1 2 DCAP8BWP7T $T=222720 427680 1 0 $X=222430 $Y=423470
X660 1 2 DCAP8BWP7T $T=226640 466880 1 0 $X=226350 $Y=462670
X661 1 2 DCAP8BWP7T $T=230000 451200 1 0 $X=229710 $Y=446990
X662 1 2 DCAP8BWP7T $T=237840 419840 0 0 $X=237550 $Y=419605
X663 1 2 DCAP8BWP7T $T=237840 459040 0 0 $X=237550 $Y=458805
X664 1 2 DCAP8BWP7T $T=238960 451200 0 0 $X=238670 $Y=450965
X665 1 2 DCAP8BWP7T $T=239520 443360 0 0 $X=239230 $Y=443125
X666 1 2 DCAP8BWP7T $T=239520 459040 1 0 $X=239230 $Y=454830
X667 1 2 DCAP8BWP7T $T=254080 427680 0 0 $X=253790 $Y=427445
X668 1 2 DCAP8BWP7T $T=256880 419840 0 0 $X=256590 $Y=419605
X669 1 2 DCAP8BWP7T $T=257440 459040 1 0 $X=257150 $Y=454830
X670 1 2 DCAP8BWP7T $T=278160 419840 0 0 $X=277870 $Y=419605
X671 1 2 DCAP8BWP7T $T=278720 459040 1 0 $X=278430 $Y=454830
X672 1 2 DCAP8BWP7T $T=279840 466880 1 0 $X=279550 $Y=462670
X673 1 2 DCAP8BWP7T $T=280960 419840 1 0 $X=280670 $Y=415630
X674 1 2 DCAP8BWP7T $T=280960 443360 1 0 $X=280670 $Y=439150
X675 1 2 DCAP8BWP7T $T=280960 451200 0 0 $X=280670 $Y=450965
X676 1 2 DCAP8BWP7T $T=280960 459040 0 0 $X=280670 $Y=458805
X677 1 2 DCAP8BWP7T $T=287120 443360 1 0 $X=286830 $Y=439150
X678 1 2 DCAP8BWP7T $T=287120 451200 0 0 $X=286830 $Y=450965
X679 1 2 DCAP8BWP7T $T=294960 419840 0 0 $X=294670 $Y=419605
X680 1 2 DCAP8BWP7T $T=302240 435520 1 0 $X=301950 $Y=431310
X681 1 2 DCAP8BWP7T $T=305040 427680 0 0 $X=304750 $Y=427445
X682 1 2 DCAP8BWP7T $T=305600 435520 0 0 $X=305310 $Y=435285
X683 1 2 DCAP8BWP7T $T=312880 419840 1 0 $X=312590 $Y=415630
X684 1 2 DCAP8BWP7T $T=319600 443360 0 0 $X=319310 $Y=443125
X685 1 2 DCAP8BWP7T $T=320720 459040 1 0 $X=320430 $Y=454830
X686 1 2 DCAP8BWP7T $T=321840 451200 0 0 $X=321550 $Y=450965
X687 1 2 DCAP8BWP7T $T=322960 435520 1 0 $X=322670 $Y=431310
X688 1 2 DCAP8BWP7T $T=323520 466880 0 0 $X=323230 $Y=466645
X689 1 2 DCAP8BWP7T $T=329120 435520 1 0 $X=328830 $Y=431310
X690 1 2 DCAP8BWP7T $T=336400 474720 1 0 $X=336110 $Y=470510
X691 1 2 DCAP8BWP7T $T=337520 435520 1 0 $X=337230 $Y=431310
X692 1 2 DCAP8BWP7T $T=346480 451200 0 0 $X=346190 $Y=450965
X693 1 2 DCAP8BWP7T $T=347040 459040 0 0 $X=346750 $Y=458805
X694 1 2 DCAP8BWP7T $T=354880 419840 1 0 $X=354590 $Y=415630
X695 1 2 DCAP8BWP7T $T=354880 443360 0 0 $X=354590 $Y=443125
X696 1 2 DCAP8BWP7T $T=362720 419840 1 0 $X=362430 $Y=415630
X697 1 2 DCAP8BWP7T $T=362720 419840 0 0 $X=362430 $Y=419605
X698 1 2 DCAP8BWP7T $T=364960 443360 0 0 $X=364670 $Y=443125
X699 1 2 DCAP8BWP7T $T=365520 451200 0 0 $X=365230 $Y=450965
X700 1 2 DCAP8BWP7T $T=371120 466880 0 0 $X=370830 $Y=466645
X701 1 2 DCAP8BWP7T $T=380080 419840 1 0 $X=379790 $Y=415630
X702 1 2 DCAP8BWP7T $T=389040 427680 0 0 $X=388750 $Y=427445
X703 1 2 DCAP8BWP7T $T=395200 443360 0 0 $X=394910 $Y=443125
X704 1 2 DCAP8BWP7T $T=396320 435520 1 0 $X=396030 $Y=431310
X705 1 2 DCAP8BWP7T $T=397440 419840 0 0 $X=397150 $Y=419605
X706 1 2 DCAP8BWP7T $T=404160 451200 1 0 $X=403870 $Y=446990
X707 1 2 DCAP8BWP7T $T=419840 443360 1 0 $X=419550 $Y=439150
X708 1 2 DCAP8BWP7T $T=426560 419840 1 0 $X=426270 $Y=415630
X709 1 2 DCAP8BWP7T $T=428800 459040 0 0 $X=428510 $Y=458805
X710 1 2 DCAP8BWP7T $T=442240 435520 0 0 $X=441950 $Y=435285
X711 1 2 DCAP8BWP7T $T=449520 427680 0 0 $X=449230 $Y=427445
X712 1 2 DCAP8BWP7T $T=449520 435520 0 0 $X=449230 $Y=435285
X713 1 2 DCAP8BWP7T $T=455120 419840 0 0 $X=454830 $Y=419605
X714 1 2 DCAP8BWP7T $T=464080 466880 1 0 $X=463790 $Y=462670
X715 2 1 DCAPBWP7T $T=22800 419840 1 0 $X=22510 $Y=415630
X716 2 1 DCAPBWP7T $T=37360 427680 0 0 $X=37070 $Y=427445
X717 2 1 DCAPBWP7T $T=45760 427680 1 0 $X=45470 $Y=423470
X718 2 1 DCAPBWP7T $T=49680 419840 1 0 $X=49390 $Y=415630
X719 2 1 DCAPBWP7T $T=49680 419840 0 0 $X=49390 $Y=419605
X720 2 1 DCAPBWP7T $T=105120 474720 1 0 $X=104830 $Y=470510
X721 2 1 DCAPBWP7T $T=121360 419840 1 0 $X=121070 $Y=415630
X722 2 1 DCAPBWP7T $T=121360 459040 1 0 $X=121070 $Y=454830
X723 2 1 DCAPBWP7T $T=125840 443360 0 0 $X=125550 $Y=443125
X724 2 1 DCAPBWP7T $T=129760 466880 1 0 $X=129470 $Y=462670
X725 2 1 DCAPBWP7T $T=131440 427680 1 0 $X=131150 $Y=423470
X726 2 1 DCAPBWP7T $T=135920 466880 1 0 $X=135630 $Y=462670
X727 2 1 DCAPBWP7T $T=140400 435520 0 0 $X=140110 $Y=435285
X728 2 1 DCAPBWP7T $T=146560 466880 0 0 $X=146270 $Y=466645
X729 2 1 DCAPBWP7T $T=158320 427680 0 0 $X=158030 $Y=427445
X730 2 1 DCAPBWP7T $T=158320 459040 1 0 $X=158030 $Y=454830
X731 2 1 DCAPBWP7T $T=174560 427680 1 0 $X=174270 $Y=423470
X732 2 1 DCAPBWP7T $T=179600 466880 0 0 $X=179310 $Y=466645
X733 2 1 DCAPBWP7T $T=180720 451200 0 0 $X=180430 $Y=450965
X734 2 1 DCAPBWP7T $T=185760 459040 0 0 $X=185470 $Y=458805
X735 2 1 DCAPBWP7T $T=200320 466880 0 0 $X=200030 $Y=466645
X736 2 1 DCAPBWP7T $T=221040 466880 1 0 $X=220750 $Y=462670
X737 2 1 DCAPBWP7T $T=222160 443360 0 0 $X=221870 $Y=443125
X738 2 1 DCAPBWP7T $T=242320 419840 0 0 $X=242030 $Y=419605
X739 2 1 DCAPBWP7T $T=242320 459040 0 0 $X=242030 $Y=458805
X740 2 1 DCAPBWP7T $T=242320 466880 1 0 $X=242030 $Y=462670
X741 2 1 DCAPBWP7T $T=247360 419840 1 0 $X=247070 $Y=415630
X742 2 1 DCAPBWP7T $T=247360 459040 0 0 $X=247070 $Y=458805
X743 2 1 DCAPBWP7T $T=249600 466880 1 0 $X=249310 $Y=462670
X744 2 1 DCAPBWP7T $T=254080 466880 0 0 $X=253790 $Y=466645
X745 2 1 DCAPBWP7T $T=266400 451200 1 0 $X=266110 $Y=446990
X746 2 1 DCAPBWP7T $T=267520 474720 1 0 $X=267230 $Y=470510
X747 2 1 DCAPBWP7T $T=284320 466880 1 0 $X=284030 $Y=462670
X748 2 1 DCAPBWP7T $T=284320 474720 1 0 $X=284030 $Y=470510
X749 2 1 DCAPBWP7T $T=296080 466880 0 0 $X=295790 $Y=466645
X750 2 1 DCAPBWP7T $T=309520 427680 0 0 $X=309230 $Y=427445
X751 2 1 DCAPBWP7T $T=326320 451200 0 0 $X=326030 $Y=450965
X752 2 1 DCAPBWP7T $T=331360 474720 1 0 $X=331070 $Y=470510
X753 2 1 DCAPBWP7T $T=333600 451200 1 0 $X=333310 $Y=446990
X754 2 1 DCAPBWP7T $T=338080 459040 1 0 $X=337790 $Y=454830
X755 2 1 DCAPBWP7T $T=340880 451200 1 0 $X=340590 $Y=446990
X756 2 1 DCAPBWP7T $T=358240 427680 0 0 $X=357950 $Y=427445
X757 2 1 DCAPBWP7T $T=359360 419840 1 0 $X=359070 $Y=415630
X758 2 1 DCAPBWP7T $T=368320 459040 0 0 $X=368030 $Y=458805
X759 2 1 DCAPBWP7T $T=373360 427680 1 0 $X=373070 $Y=423470
X760 2 1 DCAPBWP7T $T=385120 427680 1 0 $X=384830 $Y=423470
X761 2 1 DCAPBWP7T $T=389040 474720 1 0 $X=388750 $Y=470510
X762 2 1 DCAPBWP7T $T=400800 435520 1 0 $X=400510 $Y=431310
X763 2 1 DCAPBWP7T $T=410320 459040 0 0 $X=410030 $Y=458805
X764 2 1 DCAPBWP7T $T=417600 419840 1 0 $X=417310 $Y=415630
X765 2 1 DCAPBWP7T $T=432160 466880 1 0 $X=431870 $Y=462670
X766 2 1 DCAPBWP7T $T=437200 466880 0 0 $X=436910 $Y=466645
X767 2 1 DCAPBWP7T $T=464080 427680 1 0 $X=463790 $Y=423470
X768 269 265 273 271 240 266 1 2 264 AO222D0BWP7T $T=303360 427680 0 180 $X=296910 $Y=423470
X769 282 265 284 271 250 266 1 2 278 AO222D0BWP7T $T=312880 435520 0 180 $X=306430 $Y=431310
X770 298 265 290 271 256 266 1 2 286 AO222D0BWP7T $T=318480 435520 1 180 $X=312030 $Y=435285
X771 312 265 311 271 285 266 1 2 304 AO222D0BWP7T $T=338640 435520 1 180 $X=332190 $Y=435285
X772 327 265 324 271 321 266 1 2 1094 AO222D0BWP7T $T=350400 435520 0 180 $X=343950 $Y=431310
X773 323 265 326 271 315 266 1 2 1098 AO222D0BWP7T $T=348160 427680 1 0 $X=347870 $Y=423470
X774 351 265 349 271 247 266 1 2 1110 AO222D0BWP7T $T=384560 435520 1 180 $X=378110 $Y=435285
X775 354 265 350 271 263 266 1 2 1111 AO222D0BWP7T $T=385120 451200 0 180 $X=378670 $Y=446990
X776 342 265 346 271 267 266 1 2 1118 AO222D0BWP7T $T=378960 459040 1 0 $X=378670 $Y=454830
X777 364 265 361 271 287 266 1 2 1128 AO222D0BWP7T $T=395200 459040 0 0 $X=394910 $Y=458805
X778 1123 265 363 271 314 266 1 2 1129 AO222D0BWP7T $T=395760 466880 1 0 $X=395470 $Y=462670
X779 369 265 375 271 310 266 1 2 1074 AO222D0BWP7T $T=408080 443360 1 180 $X=401630 $Y=443125
X780 382 265 386 271 289 266 1 2 1141 AO222D0BWP7T $T=423200 451200 1 0 $X=422910 $Y=446990
X781 385 265 394 271 253 266 1 2 1142 AO222D0BWP7T $T=437760 419840 0 180 $X=431310 $Y=415630
X782 404 265 401 271 398 266 1 2 1146 AO222D0BWP7T $T=444480 419840 1 180 $X=438030 $Y=419605
X783 408 265 415 271 377 266 1 2 1155 AO222D0BWP7T $T=451200 451200 0 180 $X=444750 $Y=446990
X784 411 265 424 271 227 266 1 2 416 AO222D0BWP7T $T=464080 427680 0 180 $X=457630 $Y=423470
X785 412 265 421 271 249 266 1 2 1148 AO222D0BWP7T $T=464080 435520 0 180 $X=457630 $Y=431310
X786 413 265 426 271 251 266 1 2 1161 AO222D0BWP7T $T=464080 443360 0 180 $X=457630 $Y=439150
X787 431 265 423 271 374 266 1 2 1156 AO222D0BWP7T $T=464080 466880 0 180 $X=457630 $Y=462670
X788 433 265 427 271 308 266 1 2 1154 AO222D0BWP7T $T=464640 443360 1 180 $X=458190 $Y=443125
X789 420 265 428 271 283 266 1 2 1162 AO222D0BWP7T $T=465200 459040 0 180 $X=458750 $Y=454830
X790 438 265 434 271 1009 266 1 2 1164 AO222D0BWP7T $T=466320 466880 1 180 $X=459870 $Y=466645
X791 445 265 446 271 246 266 1 2 1166 AO222D0BWP7T $T=469680 459040 1 180 $X=463230 $Y=458805
X792 422 1 251 430 1165 2 1167 1168 OAI221D1BWP7T $T=461840 435520 0 0 $X=461550 $Y=435285
X793 439 265 271 429 425 266 1 2 417 AO222D1BWP7T $T=466880 419840 1 180 $X=459870 $Y=419605
X794 1 2 ICV_4 $T=44640 435520 1 0 $X=44350 $Y=431310
X795 1 2 ICV_4 $T=55840 474720 1 0 $X=55550 $Y=470510
X796 1 2 ICV_4 $T=56400 435520 0 0 $X=56110 $Y=435285
X797 1 2 ICV_4 $T=107360 427680 1 0 $X=107070 $Y=423470
X798 1 2 ICV_4 $T=145440 459040 1 0 $X=145150 $Y=454830
X799 1 2 ICV_4 $T=149360 451200 0 0 $X=149070 $Y=450965
X800 1 2 ICV_4 $T=156080 474720 1 0 $X=155790 $Y=470510
X801 1 2 ICV_4 $T=179600 435520 1 0 $X=179310 $Y=431310
X802 1 2 ICV_4 $T=223840 451200 1 0 $X=223550 $Y=446990
X803 1 2 ICV_4 $T=231120 466880 1 0 $X=230830 $Y=462670
X804 1 2 ICV_4 $T=240080 419840 1 0 $X=239790 $Y=415630
X805 1 2 ICV_4 $T=240080 427680 0 0 $X=239790 $Y=427445
X806 1 2 ICV_4 $T=249600 451200 1 0 $X=249310 $Y=446990
X807 1 2 ICV_4 $T=261360 419840 0 0 $X=261070 $Y=419605
X808 1 2 ICV_4 $T=266960 451200 0 0 $X=266670 $Y=450965
X809 1 2 ICV_4 $T=271440 443360 0 0 $X=271150 $Y=443125
X810 1 2 ICV_4 $T=274800 427680 0 0 $X=274510 $Y=427445
X811 1 2 ICV_4 $T=282080 435520 1 0 $X=281790 $Y=431310
X812 1 2 ICV_4 $T=291600 451200 1 0 $X=291310 $Y=446990
X813 1 2 ICV_4 $T=301680 443360 1 0 $X=301390 $Y=439150
X814 1 2 ICV_4 $T=324080 443360 0 0 $X=323790 $Y=443125
X815 1 2 ICV_4 $T=338080 443360 0 0 $X=337790 $Y=443125
X816 1 2 ICV_4 $T=366080 459040 1 0 $X=365790 $Y=454830
X817 1 2 ICV_4 $T=366080 466880 1 0 $X=365790 $Y=462670
X818 1 2 ICV_4 $T=366080 474720 1 0 $X=365790 $Y=470510
X819 1 2 ICV_4 $T=384560 435520 0 0 $X=384270 $Y=435285
X820 1 2 ICV_4 $T=394080 474720 1 0 $X=393790 $Y=470510
X821 1 2 ICV_4 $T=408080 419840 1 0 $X=407790 $Y=415630
X822 1 2 ICV_4 $T=408080 451200 0 0 $X=407790 $Y=450965
X823 1 2 ICV_4 $T=408080 466880 0 0 $X=407790 $Y=466645
X824 1 2 ICV_4 $T=450080 435520 1 0 $X=449790 $Y=431310
X825 1 2 ICV_4 $T=450080 459040 1 0 $X=449790 $Y=454830
X826 1 2 ICV_4 $T=450080 466880 1 0 $X=449790 $Y=462670
X827 1 2 ICV_4 $T=459600 459040 0 0 $X=459310 $Y=458805
X828 294 1080 288 2 1 1043 DFCNQD1BWP7T $T=325200 427680 0 180 $X=312590 $Y=423470
X829 294 301 288 2 1 1046 DFCNQD1BWP7T $T=325200 459040 1 180 $X=312590 $Y=458805
X830 294 1083 288 2 1 1063 DFCNQD1BWP7T $T=344800 427680 0 180 $X=332190 $Y=423470
X831 294 1094 288 2 1 262 DFCNQD1BWP7T $T=348720 419840 1 180 $X=336110 $Y=419605
X832 294 1089 288 2 1 1086 DFCNQD1BWP7T $T=349280 427680 1 180 $X=336670 $Y=427445
X833 294 1092 288 2 1 1064 DFCNQD1BWP7T $T=352080 459040 0 180 $X=339470 $Y=454830
X834 294 1079 288 2 1 1012 DFCNQD1BWP7T $T=353200 466880 0 180 $X=340590 $Y=462670
X835 294 1085 288 2 1 1069 DFCNQD1BWP7T $T=360480 466880 1 180 $X=347870 $Y=466645
X836 294 1096 288 2 1 1077 DFCNQD1BWP7T $T=366080 459040 0 180 $X=353470 $Y=454830
X837 294 1104 288 2 1 1050 DFCNQD1BWP7T $T=366080 466880 0 180 $X=353470 $Y=462670
X838 294 1106 288 2 1 1035 DFCNQD1BWP7T $T=367200 435520 0 180 $X=354590 $Y=431310
X839 294 1111 288 2 1 1107 DFCNQD1BWP7T $T=386240 459040 1 180 $X=373630 $Y=458805
X840 294 1110 288 2 1 1119 DFCNQD1BWP7T $T=378400 466880 1 0 $X=378110 $Y=462670
X841 294 1139 288 2 1 1075 DFCNQD1BWP7T $T=428240 466880 1 180 $X=415630 $Y=466645
X842 294 1138 288 2 1 1068 DFCNQD1BWP7T $T=428240 474720 0 180 $X=415630 $Y=470510
X843 294 390 288 2 1 1101 DFCNQD1BWP7T $T=430480 419840 1 180 $X=417870 $Y=419605
X844 294 1143 288 2 1 1032 DFCNQD1BWP7T $T=432160 466880 0 180 $X=419550 $Y=462670
X845 294 1144 288 2 1 1067 DFCNQD1BWP7T $T=433280 459040 0 180 $X=420670 $Y=454830
X846 294 1151 288 2 1 1017 DFCNQD1BWP7T $T=441680 451200 0 180 $X=429070 $Y=446990
X847 294 1154 288 2 1 1134 DFCNQD1BWP7T $T=447840 451200 1 180 $X=435230 $Y=450965
X848 294 1161 288 2 1 396 DFCNQD1BWP7T $T=450080 459040 0 180 $X=437470 $Y=454830
X849 294 1162 288 2 1 1130 DFCNQD1BWP7T $T=451200 466880 1 180 $X=438590 $Y=466645
X850 294 1166 288 2 1 1122 DFCNQD1BWP7T $T=470240 451200 0 180 $X=457630 $Y=446990
X851 294 1164 288 2 1 1163 DFCNQD1BWP7T $T=470800 451200 1 180 $X=458190 $Y=450965
X1100 1 2 ICV_8 $T=20000 427680 0 0 $X=19710 $Y=427445
X1101 1 2 ICV_8 $T=20000 459040 0 0 $X=19710 $Y=458805
X1102 1 2 ICV_8 $T=34000 435520 0 0 $X=33710 $Y=435285
X1103 1 2 ICV_8 $T=34000 443360 1 0 $X=33710 $Y=439150
X1104 1 2 ICV_8 $T=34000 443360 0 0 $X=33710 $Y=443125
X1105 1 2 ICV_8 $T=34000 466880 0 0 $X=33710 $Y=466645
X1106 1 2 ICV_8 $T=34000 474720 1 0 $X=33710 $Y=470510
X1107 1 2 ICV_8 $T=118000 419840 0 0 $X=117710 $Y=419605
X1108 1 2 ICV_8 $T=118000 451200 1 0 $X=117710 $Y=446990
X1109 1 2 ICV_8 $T=118000 451200 0 0 $X=117710 $Y=450965
X1110 1 2 ICV_8 $T=160000 451200 0 0 $X=159710 $Y=450965
X1111 1 2 ICV_8 $T=160000 459040 1 0 $X=159710 $Y=454830
X1112 1 2 ICV_8 $T=160000 466880 1 0 $X=159710 $Y=462670
X1113 1 2 ICV_8 $T=202000 466880 0 0 $X=201710 $Y=466645
X1114 1 2 ICV_8 $T=202000 474720 1 0 $X=201710 $Y=470510
X1115 1 2 ICV_8 $T=244000 466880 1 0 $X=243710 $Y=462670
X1116 1 2 ICV_8 $T=244000 466880 0 0 $X=243710 $Y=466645
X1117 1 2 ICV_8 $T=286000 419840 0 0 $X=285710 $Y=419605
X1118 1 2 ICV_8 $T=286000 427680 0 0 $X=285710 $Y=427445
X1119 1 2 ICV_8 $T=286000 459040 1 0 $X=285710 $Y=454830
X1120 1 2 ICV_8 $T=286000 466880 1 0 $X=285710 $Y=462670
X1121 1 2 ICV_8 $T=286000 474720 1 0 $X=285710 $Y=470510
X1122 1 2 ICV_8 $T=328000 419840 0 0 $X=327710 $Y=419605
X1123 1 2 ICV_8 $T=370000 435520 1 0 $X=369710 $Y=431310
X1124 1 2 ICV_8 $T=370000 451200 1 0 $X=369710 $Y=446990
X1125 1 2 ICV_8 $T=370000 451200 0 0 $X=369710 $Y=450965
X1126 1 2 ICV_8 $T=370000 459040 0 0 $X=369710 $Y=458805
X1127 1 2 ICV_8 $T=412000 443360 1 0 $X=411710 $Y=439150
X1128 1 2 ICV_8 $T=412000 451200 0 0 $X=411710 $Y=450965
X1129 1 2 ICV_8 $T=412000 459040 0 0 $X=411710 $Y=458805
X1130 1 2 ICV_8 $T=412000 466880 0 0 $X=411710 $Y=466645
X1131 1 2 ICV_8 $T=412000 474720 1 0 $X=411710 $Y=470510
X1132 1 2 ICV_8 $T=454000 435520 1 0 $X=453710 $Y=431310
X1133 1 2 ICV_8 $T=454000 435520 0 0 $X=453710 $Y=435285
X1134 1 2 ICV_8 $T=454000 451200 1 0 $X=453710 $Y=446990
X1135 1 2 ICV_8 $T=454000 466880 1 0 $X=453710 $Y=462670
X1136 1 2 ICV_9 $T=34000 451200 1 0 $X=33710 $Y=446990
X1137 1 2 ICV_9 $T=34000 459040 1 0 $X=33710 $Y=454830
X1138 1 2 ICV_9 $T=34000 459040 0 0 $X=33710 $Y=458805
X1139 1 2 ICV_9 $T=34000 466880 1 0 $X=33710 $Y=462670
X1140 1 2 ICV_9 $T=160000 459040 0 0 $X=159710 $Y=458805
X1141 1 2 ICV_9 $T=160000 474720 1 0 $X=159710 $Y=470510
X1142 1 2 ICV_9 $T=202000 435520 1 0 $X=201710 $Y=431310
X1143 1 2 ICV_9 $T=244000 427680 1 0 $X=243710 $Y=423470
X1144 1 2 ICV_9 $T=244000 427680 0 0 $X=243710 $Y=427445
X1145 1 2 ICV_9 $T=244000 435520 1 0 $X=243710 $Y=431310
X1146 1 2 ICV_9 $T=244000 435520 0 0 $X=243710 $Y=435285
X1147 1 2 ICV_9 $T=244000 451200 1 0 $X=243710 $Y=446990
X1148 1 2 ICV_9 $T=244000 459040 1 0 $X=243710 $Y=454830
X1149 1 2 ICV_9 $T=286000 435520 0 0 $X=285710 $Y=435285
X1150 1 2 ICV_9 $T=286000 443360 0 0 $X=285710 $Y=443125
X1151 1 2 ICV_9 $T=286000 451200 1 0 $X=285710 $Y=446990
X1152 1 2 ICV_9 $T=328000 419840 1 0 $X=327710 $Y=415630
X1153 1 2 ICV_9 $T=328000 427680 0 0 $X=327710 $Y=427445
X1154 1 2 ICV_9 $T=328000 443360 1 0 $X=327710 $Y=439150
X1155 1 2 ICV_9 $T=328000 451200 1 0 $X=327710 $Y=446990
X1156 1 2 ICV_9 $T=328000 451200 0 0 $X=327710 $Y=450965
X1157 1 2 ICV_9 $T=328000 459040 0 0 $X=327710 $Y=458805
X1158 1 2 ICV_9 $T=328000 466880 1 0 $X=327710 $Y=462670
X1159 1 2 ICV_9 $T=328000 466880 0 0 $X=327710 $Y=466645
X1160 1 2 ICV_9 $T=370000 443360 1 0 $X=369710 $Y=439150
X1161 1 2 ICV_9 $T=370000 459040 1 0 $X=369710 $Y=454830
X1162 1 2 ICV_9 $T=370000 466880 1 0 $X=369710 $Y=462670
X1163 1 2 ICV_9 $T=370000 474720 1 0 $X=369710 $Y=470510
X1164 1 2 ICV_9 $T=412000 419840 1 0 $X=411710 $Y=415630
X1165 1 2 ICV_9 $T=412000 419840 0 0 $X=411710 $Y=419605
X1166 1 2 ICV_9 $T=412000 435520 0 0 $X=411710 $Y=435285
X1167 1 2 ICV_9 $T=412000 443360 0 0 $X=411710 $Y=443125
X1168 1 2 ICV_9 $T=412000 459040 1 0 $X=411710 $Y=454830
X1169 1 2 ICV_9 $T=412000 466880 1 0 $X=411710 $Y=462670
X1170 1 2 ICV_9 $T=454000 427680 0 0 $X=453710 $Y=427445
X1171 1 2 ICV_9 $T=454000 459040 0 0 $X=453710 $Y=458805
X1172 1 2 ICV_10 $T=20000 451200 1 0 $X=19710 $Y=446990
X1173 1 2 ICV_10 $T=20000 466880 1 0 $X=19710 $Y=462670
X1174 1 2 ICV_10 $T=34000 419840 1 0 $X=33710 $Y=415630
X1175 1 2 ICV_10 $T=34000 427680 0 0 $X=33710 $Y=427445
X1176 1 2 ICV_10 $T=34000 451200 0 0 $X=33710 $Y=450965
X1177 1 2 ICV_10 $T=118000 419840 1 0 $X=117710 $Y=415630
X1178 1 2 ICV_10 $T=118000 427680 0 0 $X=117710 $Y=427445
X1179 1 2 ICV_10 $T=118000 459040 1 0 $X=117710 $Y=454830
X1180 1 2 ICV_10 $T=118000 466880 0 0 $X=117710 $Y=466645
X1181 1 2 ICV_10 $T=118000 474720 1 0 $X=117710 $Y=470510
X1182 1 2 ICV_10 $T=160000 443360 0 0 $X=159710 $Y=443125
X1183 1 2 ICV_10 $T=202000 435520 0 0 $X=201710 $Y=435285
X1184 1 2 ICV_10 $T=202000 459040 1 0 $X=201710 $Y=454830
X1185 1 2 ICV_10 $T=244000 419840 1 0 $X=243710 $Y=415630
X1186 1 2 ICV_10 $T=244000 443360 0 0 $X=243710 $Y=443125
X1187 1 2 ICV_10 $T=244000 459040 0 0 $X=243710 $Y=458805
X1188 1 2 ICV_10 $T=286000 427680 1 0 $X=285710 $Y=423470
X1189 1 2 ICV_10 $T=328000 427680 1 0 $X=327710 $Y=423470
X1190 1 2 ICV_10 $T=328000 435520 0 0 $X=327710 $Y=435285
X1191 1 2 ICV_10 $T=328000 474720 1 0 $X=327710 $Y=470510
X1192 1 2 ICV_10 $T=370000 427680 1 0 $X=369710 $Y=423470
X1193 1 2 ICV_10 $T=412000 451200 1 0 $X=411710 $Y=446990
X1194 1 2 ICV_10 $T=454000 459040 1 0 $X=453710 $Y=454830
X1236 1 2 ICV_13 $T=30640 427680 0 0 $X=30350 $Y=427445
X1237 1 2 ICV_13 $T=30640 443360 1 0 $X=30350 $Y=439150
X1238 1 2 ICV_13 $T=30640 451200 0 0 $X=30350 $Y=450965
X1239 1 2 ICV_13 $T=46320 466880 1 0 $X=46030 $Y=462670
X1240 1 2 ICV_13 $T=50800 466880 0 0 $X=50510 $Y=466645
X1241 1 2 ICV_13 $T=114640 451200 1 0 $X=114350 $Y=446990
X1242 1 2 ICV_13 $T=119120 443360 0 0 $X=118830 $Y=443125
X1243 1 2 ICV_13 $T=132000 419840 0 0 $X=131710 $Y=419605
X1244 1 2 ICV_13 $T=133120 435520 0 0 $X=132830 $Y=435285
X1245 1 2 ICV_13 $T=141520 451200 0 0 $X=141230 $Y=450965
X1246 1 2 ICV_13 $T=142640 459040 0 0 $X=142350 $Y=458805
X1247 1 2 ICV_13 $T=156640 435520 0 0 $X=156350 $Y=435285
X1248 1 2 ICV_13 $T=161120 435520 1 0 $X=160830 $Y=431310
X1249 1 2 ICV_13 $T=230000 459040 1 0 $X=229710 $Y=454830
X1250 1 2 ICV_13 $T=240640 427680 1 0 $X=240350 $Y=423470
X1251 1 2 ICV_13 $T=261920 459040 1 0 $X=261630 $Y=454830
X1252 1 2 ICV_13 $T=282640 419840 0 0 $X=282350 $Y=419605
X1253 1 2 ICV_13 $T=291600 443360 0 0 $X=291310 $Y=443125
X1254 1 2 ICV_13 $T=333600 427680 0 0 $X=333310 $Y=427445
X1255 1 2 ICV_13 $T=333600 466880 0 0 $X=333310 $Y=466645
X1256 1 2 ICV_13 $T=338640 419840 1 0 $X=338350 $Y=415630
X1257 1 2 ICV_13 $T=344800 427680 1 0 $X=344510 $Y=423470
X1258 1 2 ICV_13 $T=350960 451200 0 0 $X=350670 $Y=450965
X1259 1 2 ICV_13 $T=357680 427680 1 0 $X=357390 $Y=423470
X1260 1 2 ICV_13 $T=359360 451200 0 0 $X=359070 $Y=450965
X1261 1 2 ICV_13 $T=382880 474720 1 0 $X=382590 $Y=470510
X1262 1 2 ICV_13 $T=408640 443360 1 0 $X=408350 $Y=439150
X1263 1 2 ICV_13 $T=408640 443360 0 0 $X=408350 $Y=443125
X1264 1 2 ICV_13 $T=408640 451200 1 0 $X=408350 $Y=446990
X1265 1 2 ICV_13 $T=417600 459040 1 0 $X=417310 $Y=454830
X1266 1 2 ICV_13 $T=420960 419840 1 0 $X=420670 $Y=415630
X1267 1 2 ICV_13 $T=441680 451200 1 0 $X=441390 $Y=446990
X1268 1 2 ICV_13 $T=450640 443360 0 0 $X=450350 $Y=443125
X1269 786 232 2 232 1004 786 1 MAOI22D1BWP7T $T=249600 427680 0 0 $X=249310 $Y=427445
X1270 1006 963 2 963 242 1006 1 MAOI22D1BWP7T $T=253520 419840 1 0 $X=253230 $Y=415630
X1271 908 987 2 987 1016 908 1 MAOI22D1BWP7T $T=255760 466880 0 0 $X=255470 $Y=466645
X1272 224 958 2 958 1026 224 1 MAOI22D1BWP7T $T=267520 443360 0 180 $X=262750 $Y=439150
X1273 364 362 2 364 1097 362 1 MAOI22D1BWP7T $T=401920 443360 0 180 $X=397150 $Y=439150
X1274 1127 367 2 367 1099 1127 1 MAOI22D1BWP7T $T=404160 435520 1 180 $X=399390 $Y=435285
X1275 368 371 2 371 1078 368 1 MAOI22D1BWP7T $T=406400 419840 1 180 $X=401630 $Y=419605
X1276 327 373 2 327 1093 373 1 MAOI22D1BWP7T $T=409200 435520 0 180 $X=404430 $Y=431310
X1277 1136 382 2 382 1116 1136 1 MAOI22D1BWP7T $T=422640 443360 1 180 $X=417870 $Y=443125
X1278 412 407 2 412 1114 407 1 MAOI22D1BWP7T $T=451200 427680 0 180 $X=446430 $Y=423470
X1279 1051 261 1 259 257 2 IOA21D0BWP7T $T=294400 419840 0 180 $X=290750 $Y=415630
X1280 1055 265 1 268 1057 2 IOA21D0BWP7T $T=297200 419840 1 0 $X=296910 $Y=415630
X1281 1081 265 1 1076 293 2 IOA21D0BWP7T $T=322960 435520 0 180 $X=319310 $Y=431310
X1282 1082 265 1 1079 300 2 IOA21D0BWP7T $T=324640 435520 1 180 $X=320990 $Y=435285
X1283 1088 265 1 1085 307 2 IOA21D0BWP7T $T=338640 451200 0 180 $X=334990 $Y=446990
X1284 1093 265 1 1089 317 2 IOA21D0BWP7T $T=344240 435520 1 180 $X=340590 $Y=435285
X1285 1095 265 1 1092 1090 2 IOA21D0BWP7T $T=345920 451200 0 180 $X=342270 $Y=446990
X1286 1097 265 1 1096 325 2 IOA21D0BWP7T $T=352080 451200 0 180 $X=348430 $Y=446990
X1287 1112 265 1 1106 344 2 IOA21D0BWP7T $T=380640 435520 0 180 $X=376990 $Y=431310
X1288 1114 265 1 1080 347 2 IOA21D0BWP7T $T=385120 427680 0 180 $X=381470 $Y=423470
X1289 1124 265 1 1115 1120 2 IOA21D0BWP7T $T=395200 443360 1 180 $X=391550 $Y=443125
X1290 1137 265 1 1135 380 2 IOA21D0BWP7T $T=419840 451200 0 180 $X=416190 $Y=446990
X1291 1145 265 1 1139 391 2 IOA21D0BWP7T $T=431040 443360 0 180 $X=427390 $Y=439150
X1292 1149 265 1 1144 1140 2 IOA21D0BWP7T $T=437200 443360 0 180 $X=433550 $Y=439150
X1293 1152 265 1 1151 397 2 IOA21D0BWP7T $T=442240 435520 1 180 $X=438590 $Y=435285
X1294 1157 265 1 1143 399 2 IOA21D0BWP7T $T=444480 443360 0 180 $X=440830 $Y=439150
X1295 1158 265 1 1153 1150 2 IOA21D0BWP7T $T=446160 435520 0 180 $X=442510 $Y=431310
X1296 1159 265 1 1131 402 2 IOA21D0BWP7T $T=446720 419840 0 180 $X=443070 $Y=415630
X1297 1160 265 1 1138 403 2 IOA21D0BWP7T $T=446720 427680 0 180 $X=443070 $Y=423470
X1298 7 1 2 4 INVD1BWP7T $T=22800 419840 0 180 $X=20830 $Y=415630
X1299 480 1 2 458 INVD1BWP7T $T=28960 443360 1 180 $X=26990 $Y=443125
X1300 3 1 2 19 INVD1BWP7T $T=28960 435520 0 0 $X=28670 $Y=435285
X1301 493 1 2 476 INVD1BWP7T $T=39600 443360 0 180 $X=37630 $Y=439150
X1302 497 1 2 496 INVD1BWP7T $T=42960 435520 1 0 $X=42670 $Y=431310
X1303 503 1 2 519 INVD1BWP7T $T=48560 435520 1 0 $X=48270 $Y=431310
X1304 35 1 2 510 INVD1BWP7T $T=54160 459040 0 180 $X=52190 $Y=454830
X1305 531 1 2 524 INVD1BWP7T $T=56400 466880 1 0 $X=56110 $Y=462670
X1306 549 1 2 501 INVD1BWP7T $T=59200 451200 1 180 $X=57230 $Y=450965
X1307 44 1 2 569 INVD1BWP7T $T=62000 443360 0 0 $X=61710 $Y=443125
X1308 614 1 2 616 INVD1BWP7T $T=83840 459040 0 0 $X=83550 $Y=458805
X1309 65 1 2 606 INVD1BWP7T $T=100080 427680 0 0 $X=99790 $Y=427445
X1310 633 1 2 690 INVD1BWP7T $T=105120 427680 0 0 $X=104830 $Y=427445
X1311 559 1 2 638 INVD1BWP7T $T=105120 435520 0 0 $X=104830 $Y=435285
X1312 731 1 2 512 INVD1BWP7T $T=125840 419840 1 180 $X=123870 $Y=419605
X1313 687 1 2 735 INVD1BWP7T $T=135360 451200 0 0 $X=135070 $Y=450965
X1314 744 1 2 677 INVD1BWP7T $T=138160 466880 1 180 $X=136190 $Y=466645
X1315 105 1 2 768 INVD1BWP7T $T=147680 459040 1 180 $X=145710 $Y=458805
X1316 132 1 2 112 INVD1BWP7T $T=157200 419840 0 180 $X=155230 $Y=415630
X1317 129 1 2 808 INVD1BWP7T $T=163920 459040 1 0 $X=163630 $Y=454830
X1318 131 1 2 809 INVD1BWP7T $T=165040 443360 0 0 $X=164750 $Y=443125
X1319 142 1 2 145 INVD1BWP7T $T=167280 435520 0 0 $X=166990 $Y=435285
X1320 157 1 2 827 INVD1BWP7T $T=175120 451200 0 180 $X=173150 $Y=446990
X1321 161 1 2 860 INVD1BWP7T $T=179600 427680 0 0 $X=179310 $Y=427445
X1322 169 1 2 784 INVD1BWP7T $T=185200 435520 0 180 $X=183230 $Y=431310
X1323 895 1 2 884 INVD1BWP7T $T=207600 466880 0 180 $X=205630 $Y=462670
X1324 936 1 2 915 INVD1BWP7T $T=212640 451200 0 0 $X=212350 $Y=450965
X1325 949 1 2 880 INVD1BWP7T $T=216000 451200 1 180 $X=214030 $Y=450965
X1326 965 1 2 978 INVD1BWP7T $T=226640 435520 1 0 $X=226350 $Y=431310
X1327 221 1 2 975 INVD1BWP7T $T=230000 459040 0 180 $X=228030 $Y=454830
X1328 89 1 2 219 INVD1BWP7T $T=231680 435520 0 180 $X=229710 $Y=431310
X1329 92 1 2 980 INVD1BWP7T $T=231680 451200 1 180 $X=229710 $Y=450965
X1330 220 1 2 987 INVD1BWP7T $T=236720 443360 1 0 $X=236430 $Y=439150
X1331 291 1 2 1073 INVD1BWP7T $T=317360 451200 1 0 $X=317070 $Y=446990
X1332 342 1 2 340 INVD1BWP7T $T=376720 427680 0 180 $X=374750 $Y=423470
X1333 400 1 2 1136 INVD1BWP7T $T=440560 427680 1 180 $X=438590 $Y=427445
X1334 1 2 ICV_14 $T=133680 427680 0 0 $X=133390 $Y=427445
X1335 1 2 ICV_14 $T=143760 435520 1 0 $X=143470 $Y=431310
X1336 1 2 ICV_14 $T=217680 474720 1 0 $X=217390 $Y=470510
X1337 1 2 ICV_14 $T=238400 435520 1 0 $X=238110 $Y=431310
X1338 1 2 ICV_14 $T=238400 435520 0 0 $X=238110 $Y=435285
X1339 1 2 ICV_14 $T=238400 443360 1 0 $X=238110 $Y=439150
X1340 1 2 ICV_14 $T=262480 459040 0 0 $X=262190 $Y=458805
X1341 1 2 ICV_14 $T=264160 427680 1 0 $X=263870 $Y=423470
X1342 1 2 ICV_14 $T=280400 427680 0 0 $X=280110 $Y=427445
X1343 1 2 ICV_14 $T=280400 435520 0 0 $X=280110 $Y=435285
X1344 1 2 ICV_14 $T=280400 443360 0 0 $X=280110 $Y=443125
X1345 1 2 ICV_14 $T=303360 419840 1 0 $X=303070 $Y=415630
X1346 1 2 ICV_14 $T=303360 419840 0 0 $X=303070 $Y=419605
X1347 1 2 ICV_14 $T=322400 419840 1 0 $X=322110 $Y=415630
X1348 1 2 ICV_14 $T=364400 427680 1 0 $X=364110 $Y=423470
X1349 1 2 ICV_14 $T=387360 435520 1 0 $X=387070 $Y=431310
X1350 1 2 ICV_14 $T=398000 427680 1 0 $X=397710 $Y=423470
X1351 1 2 ICV_14 $T=406400 419840 0 0 $X=406110 $Y=419605
X1352 1 2 ICV_14 $T=433280 435520 0 0 $X=432990 $Y=435285
X1353 1 2 ICV_14 $T=437200 435520 1 0 $X=436910 $Y=431310
X1354 1 2 ICV_14 $T=437760 419840 1 0 $X=437470 $Y=415630
X1355 1 2 294 292 288 1066 ICV_15 $T=320720 466880 0 180 $X=308110 $Y=462670
X1356 1 2 294 1074 288 280 ICV_15 $T=321280 419840 1 180 $X=308670 $Y=419605
X1357 1 2 294 1076 288 1042 ICV_15 $T=323520 427680 1 180 $X=310910 $Y=427445
X1358 1 2 294 1100 288 1061 ICV_15 $T=363840 459040 1 180 $X=351230 $Y=458805
X1359 1 2 294 1103 288 1060 ICV_15 $T=365520 435520 1 180 $X=352910 $Y=435285
X1360 1 2 294 1113 288 1072 ICV_15 $T=386240 451200 1 180 $X=373630 $Y=450965
X1361 1 2 294 1115 288 1091 ICV_15 $T=387360 443360 1 180 $X=374750 $Y=443125
X1362 1 2 294 1118 288 1109 ICV_15 $T=390720 466880 1 180 $X=378110 $Y=466645
X1363 1 2 294 1129 288 355 ICV_15 $T=403600 451200 1 180 $X=390990 $Y=450965
X1364 1 2 294 1131 288 1002 ICV_15 $T=404720 459040 0 180 $X=392110 $Y=454830
X1365 1 2 294 1135 288 1019 ICV_15 $T=428240 451200 1 180 $X=415630 $Y=450965
X1366 1 2 294 1142 288 1125 ICV_15 $T=432160 427680 1 180 $X=419550 $Y=427445
X1367 1 2 294 1146 336 1133 ICV_15 $T=434960 427680 0 180 $X=422350 $Y=423470
X1368 1 2 294 1153 288 1070 ICV_15 $T=446160 443360 1 180 $X=433550 $Y=443125
X1369 1 2 294 1155 288 1147 ICV_15 $T=447280 459040 1 180 $X=434670 $Y=458805
X1370 1 2 294 1156 288 1132 ICV_15 $T=447280 474720 0 180 $X=434670 $Y=470510
X1371 393 302 1 2 BUFFD10BWP7T $T=433840 466880 1 0 $X=433550 $Y=462670
X1372 222 217 1 2 BUFFD2BWP7T $T=226640 474720 0 180 $X=222990 $Y=470510
X1373 1030 308 1 2 BUFFD2BWP7T $T=333040 474720 1 0 $X=332750 $Y=470510
X1374 1056 310 1 2 BUFFD2BWP7T $T=334720 459040 0 0 $X=334430 $Y=458805
X1375 1101 332 1 2 BUFFD2BWP7T $T=362720 419840 1 180 $X=359070 $Y=419605
X1376 1122 296 1 2 BUFFD2BWP7T $T=394080 474720 0 180 $X=390430 $Y=470510
X1377 1125 331 1 2 BUFFD2BWP7T $T=396320 435520 0 180 $X=392670 $Y=431310
X1378 1065 374 1 2 BUFFD2BWP7T $T=402480 474720 1 0 $X=402190 $Y=470510
X1379 1133 372 1 2 BUFFD2BWP7T $T=406960 427680 0 180 $X=403310 $Y=423470
X1380 1071 377 1 2 BUFFD2BWP7T $T=405840 474720 1 0 $X=405550 $Y=470510
X1381 1147 392 1 2 BUFFD2BWP7T $T=432720 466880 1 180 $X=429070 $Y=466645
X1382 294 1098 288 318 1 2 DFCNQD2BWP7T $T=354880 419840 0 180 $X=341710 $Y=415630
X1383 294 359 288 322 1 2 DFCNQD2BWP7T $T=399120 419840 0 180 $X=385950 $Y=415630
X1384 294 1128 288 356 1 2 DFCNQD2BWP7T $T=404160 451200 0 180 $X=390990 $Y=446990
X1385 294 1141 288 384 1 2 DFCNQD2BWP7T $T=433280 435520 1 180 $X=420110 $Y=435285
X1386 294 1148 336 389 1 2 DFCNQD2BWP7T $T=437200 435520 0 180 $X=424030 $Y=431310
X1387 1 2 DCAP16BWP7T $T=214880 451200 1 0 $X=214590 $Y=446990
X1388 1 2 DCAP16BWP7T $T=245120 419840 0 0 $X=244830 $Y=419605
X1389 1 2 DCAP16BWP7T $T=258000 419840 1 0 $X=257710 $Y=415630
X1390 1 2 DCAP16BWP7T $T=262480 443360 0 0 $X=262190 $Y=443125
X1391 1 2 DCAP16BWP7T $T=272000 419840 1 0 $X=271710 $Y=415630
X1392 1 2 DCAP16BWP7T $T=287120 459040 0 0 $X=286830 $Y=458805
X1393 1 2 DCAP16BWP7T $T=287120 466880 0 0 $X=286830 $Y=466645
X1394 1 2 DCAP16BWP7T $T=296080 427680 0 0 $X=295790 $Y=427445
X1395 1 2 DCAP16BWP7T $T=303360 427680 1 0 $X=303070 $Y=423470
X1396 1 2 DCAP16BWP7T $T=308400 451200 1 0 $X=308110 $Y=446990
X1397 1 2 DCAP16BWP7T $T=319040 443360 1 0 $X=318750 $Y=439150
X1398 1 2 DCAP16BWP7T $T=319040 451200 1 0 $X=318750 $Y=446990
X1399 1 2 DCAP16BWP7T $T=329120 443360 0 0 $X=328830 $Y=443125
X1400 1 2 DCAP16BWP7T $T=329120 459040 1 0 $X=328830 $Y=454830
X1401 1 2 DCAP16BWP7T $T=338080 459040 0 0 $X=337790 $Y=458805
X1402 1 2 DCAP16BWP7T $T=348720 419840 0 0 $X=348430 $Y=419605
X1403 1 2 DCAP16BWP7T $T=349280 427680 0 0 $X=348990 $Y=427445
X1404 1 2 DCAP16BWP7T $T=350400 474720 1 0 $X=350110 $Y=470510
X1405 1 2 DCAP16BWP7T $T=359920 443360 1 0 $X=359630 $Y=439150
X1406 1 2 DCAP16BWP7T $T=360480 466880 0 0 $X=360190 $Y=466645
X1407 1 2 DCAP16BWP7T $T=371120 419840 1 0 $X=370830 $Y=415630
X1408 1 2 DCAP16BWP7T $T=371120 427680 0 0 $X=370830 $Y=427445
X1409 1 2 DCAP16BWP7T $T=379520 419840 0 0 $X=379230 $Y=419605
X1410 1 2 DCAP16BWP7T $T=385680 443360 1 0 $X=385390 $Y=439150
X1411 1 2 DCAP16BWP7T $T=386240 459040 0 0 $X=385950 $Y=458805
X1412 1 2 DCAP16BWP7T $T=389040 427680 1 0 $X=388750 $Y=423470
X1413 1 2 DCAP16BWP7T $T=399120 419840 1 0 $X=398830 $Y=415630
X1414 1 2 DCAP16BWP7T $T=401360 459040 0 0 $X=401070 $Y=458805
X1415 1 2 DCAP16BWP7T $T=401920 466880 1 0 $X=401630 $Y=462670
X1416 1 2 DCAP16BWP7T $T=413120 435520 1 0 $X=412830 $Y=431310
X1417 1 2 DCAP16BWP7T $T=419840 459040 0 0 $X=419550 $Y=458805
X1418 494 1 2 505 CKND1BWP7T $T=42960 451200 1 0 $X=42670 $Y=446990
X1419 460 1 2 508 CKND1BWP7T $T=43520 435520 0 0 $X=43230 $Y=435285
X1420 75 1 2 601 CKND1BWP7T $T=102320 443360 1 180 $X=100350 $Y=443125
X1421 84 1 2 86 CKND1BWP7T $T=128640 419840 0 180 $X=126670 $Y=415630
X1422 80 1 2 728 CKND1BWP7T $T=127520 419840 0 0 $X=127230 $Y=419605
X1423 758 1 2 722 CKND1BWP7T $T=138160 435520 1 180 $X=136190 $Y=435285
X1424 756 1 2 100 CKND1BWP7T $T=143760 443360 0 0 $X=143470 $Y=443125
X1425 98 1 2 782 CKND1BWP7T $T=147680 443360 1 0 $X=147390 $Y=439150
X1426 216 1 2 970 CKND1BWP7T $T=222720 466880 1 0 $X=222430 $Y=462670
X1427 723 1 2 982 CKND1BWP7T $T=236160 459040 0 0 $X=235870 $Y=458805
X1428 236 1 2 998 CKND1BWP7T $T=249600 459040 1 0 $X=249310 $Y=454830
X1429 786 1 2 237 CKND1BWP7T $T=253520 435520 1 0 $X=253230 $Y=431310
X1430 241 1 2 1006 CKND1BWP7T $T=256880 419840 1 180 $X=254910 $Y=419605
X1431 383 1 2 1126 CKND1BWP7T $T=420960 419840 0 180 $X=418990 $Y=415630
X1432 378 381 1 2 INVD4BWP7T $T=415920 459040 0 0 $X=415630 $Y=458805
X1433 1109 1 2 339 BUFFD3BWP7T $T=377840 451200 0 180 $X=373630 $Y=446990
X1434 1130 1 2 366 BUFFD3BWP7T $T=401920 474720 0 180 $X=397710 $Y=470510
X1435 1132 365 1 2 BUFFD12BWP7T $T=408080 466880 1 180 $X=395470 $Y=466645
X1436 366 1126 742 1 2 CKXOR2D4BWP7T $T=407520 427680 1 180 $X=394910 $Y=427445
X1437 216 221 2 970 1 975 977 AOI22D1BWP7T $T=225520 459040 0 0 $X=225230 $Y=458805
X1438 972 220 2 984 1 987 233 AOI22D1BWP7T $T=232800 443360 1 0 $X=232510 $Y=439150
X1439 999 982 2 235 1 723 1001 AOI22D1BWP7T $T=247920 466880 0 0 $X=247630 $Y=466645
X1440 981 998 2 771 1 236 1000 AOI22D1BWP7T $T=253520 459040 1 0 $X=253230 $Y=454830
X1441 235 1024 2 999 1 908 1028 AOI22D1BWP7T $T=263600 474720 1 0 $X=263310 $Y=470510
X1442 786 973 2 237 1 1020 1038 AOI22D1BWP7T $T=268080 435520 0 0 $X=267790 $Y=435285
X1443 266 322 2 271 1 320 1090 AOI22D1BWP7T $T=349280 443360 0 180 $X=345070 $Y=439150
X1444 266 357 2 271 1 1121 1120 AOI22D1BWP7T $T=395200 419840 1 180 $X=390990 $Y=419605
X1445 297 1099 2 333 1104 1 OAI21D1BWP7T $T=363280 427680 1 180 $X=359630 $Y=427445
X1446 297 1102 2 1105 1100 1 OAI21D1BWP7T $T=361040 427680 1 0 $X=360750 $Y=423470
X1447 297 1116 2 1117 1113 1 OAI21D1BWP7T $T=384000 435520 1 0 $X=383710 $Y=431310
X1448 28 2 294 1 CKND12BWP7T $T=380080 427680 0 0 $X=379790 $Y=427445
X1449 302 288 1 2 BUFFD8BWP7T $T=325200 474720 0 180 $X=315950 $Y=470510
X1450 316 348 1 2 BUFFD8BWP7T $T=376720 443360 1 0 $X=376430 $Y=439150
X1451 271 2 265 316 1 NR2D4BWP7T $T=382880 474720 0 180 $X=375870 $Y=470510
X1452 907 896 934 1 2 957 AO21D0BWP7T $T=214880 443360 1 0 $X=214590 $Y=439150
X1453 265 1108 341 1 2 1103 AO21D0BWP7T $T=377280 435520 0 180 $X=373630 $Y=431310
X1454 319 265 1 2 BUFFD6BWP7T $T=343680 474720 1 0 $X=343390 $Y=470510
X1455 302 336 1 2 BUFFD6BWP7T $T=366080 474720 0 180 $X=359070 $Y=470510
X1456 464 8 2 1 INVD2BWP7T $T=24480 435520 0 180 $X=21950 $Y=431310
X1457 137 843 2 1 INVD2BWP7T $T=191360 427680 0 0 $X=191070 $Y=427445
X1458 234 229 2 1 INVD2BWP7T $T=251280 419840 0 180 $X=248750 $Y=415630
X1459 771 981 2 1 INVD2BWP7T $T=251840 435520 0 180 $X=249310 $Y=431310
X1460 265 297 2 1 INVD2BWP7T $T=357680 427680 0 180 $X=355150 $Y=423470
X1461 963 232 1 2 230 CKXOR2D1BWP7T $T=240080 419840 0 180 $X=234750 $Y=415630
X1462 755 991 1 2 996 CKXOR2D1BWP7T $T=235040 466880 1 0 $X=234750 $Y=462670
X1463 92 100 1 2 997 CKXOR2D1BWP7T $T=236160 474720 1 0 $X=235870 $Y=470510
X1464 296 1073 1 2 954 CKXOR2D1BWP7T $T=320720 459040 0 180 $X=315390 $Y=454830
X1465 330 329 1 2 964 CKXOR2D1BWP7T $T=359360 451200 1 180 $X=354030 $Y=450965
X1466 331 328 757 1 2 CKXOR2D2BWP7T $T=359920 443360 0 180 $X=353470 $Y=439150
X1467 2 1 DCAP32BWP7T $T=245120 443360 1 0 $X=244830 $Y=439150
X1468 2 1 DCAP32BWP7T $T=352080 451200 1 0 $X=351790 $Y=446990
X1469 219 224 983 218 981 1 2 XNR4D1BWP7T $T=225520 435520 0 0 $X=225230 $Y=435285
X1470 780 1091 314 1053 1044 1 2 XNR4D1BWP7T $T=346480 451200 1 180 $X=333310 $Y=450965
X1471 969 1086 321 1053 218 1 2 XNR4D1BWP7T $T=342000 443360 0 0 $X=341710 $Y=443125
X1472 316 1 2 266 BUFFD5BWP7T $T=339760 466880 0 180 $X=333310 $Y=462670
X1473 602 718 553 608 1 2 OAI21D0BWP7T $T=107920 466880 0 0 $X=107630 $Y=466645
X1474 744 760 740 720 1 2 OAI21D0BWP7T $T=139840 459040 0 180 $X=136750 $Y=454830
X1475 1078 299 297 295 1 2 OAI21D0BWP7T $T=322400 419840 0 180 $X=319310 $Y=415630
X1476 1084 1083 297 303 1 2 OAI21D0BWP7T $T=334720 419840 1 180 $X=331630 $Y=419605
X1477 1018 1012 1003 218 100 1 2 XNR4D0BWP7T $T=260800 474720 0 180 $X=247630 $Y=470510
X1478 1007 238 1021 245 1016 1 2 XNR4D0BWP7T $T=253520 451200 1 0 $X=253230 $Y=446990
X1479 238 1003 1023 1016 1011 1 2 XNR4D0BWP7T $T=254080 451200 0 0 $X=253790 $Y=450965
X1480 1015 979 1030 995 997 1 2 XNR4D0BWP7T $T=260240 466880 0 0 $X=259950 $Y=466645
X1481 242 1031 1034 1042 974 1 2 XNR4D0BWP7T $T=265280 419840 0 0 $X=264990 $Y=419605
X1482 1000 1032 1036 243 218 1 2 XNR4D0BWP7T $T=266960 466880 1 0 $X=266670 $Y=462670
X1483 1046 979 1040 248 995 1 2 XNR4D0BWP7T $T=280960 459040 1 180 $X=267790 $Y=458805
X1484 1049 1050 1056 977 996 1 2 XNR4D0BWP7T $T=289920 466880 1 0 $X=289630 $Y=462670
X1485 1061 243 1052 235 958 1 2 XNR4D0BWP7T $T=302800 474720 0 180 $X=289630 $Y=470510
X1486 1059 1064 1058 1039 248 1 2 XNR4D0BWP7T $T=308400 451200 0 180 $X=295230 $Y=446990
X1487 1018 992 1065 1001 1068 1 2 XNR4D0BWP7T $T=297760 466880 0 0 $X=297470 $Y=466645
X1488 996 1067 1062 1011 218 1 2 XNR4D0BWP7T $T=312880 459040 0 180 $X=299710 $Y=454830
X1489 983 1075 1071 975 1048 1 2 XNR4D0BWP7T $T=323520 466880 1 180 $X=310350 $Y=466645
X1490 993 989 227 978 963 1 2 XNR4D2BWP7T $T=240080 427680 1 180 $X=226350 $Y=427445
X1491 1026 1017 1009 985 234 1 2 XNR4D2BWP7T $T=263600 435520 1 180 $X=249870 $Y=435285
X1492 967 244 240 985 981 1 2 XNR4D2BWP7T $T=264160 427680 0 180 $X=250430 $Y=423470
X1493 1004 967 247 1035 241 1 2 XNR4D2BWP7T $T=261360 427680 0 0 $X=261070 $Y=427445
X1494 1021 780 250 975 230 1 2 XNR4D2BWP7T $T=265280 459040 1 0 $X=264990 $Y=454830
X1495 973 1036 251 252 990 1 2 XNR4D2BWP7T $T=267520 443360 1 0 $X=267230 $Y=439150
X1496 974 1043 249 1039 1020 1 2 XNR4D2BWP7T $T=282080 435520 0 180 $X=268350 $Y=431310
X1497 1029 989 253 254 1047 1 2 XNR4D2BWP7T $T=269760 427680 1 0 $X=269470 $Y=423470
X1498 1029 1054 272 780 1063 1 2 XNR4D2BWP7T $T=292160 435520 0 0 $X=291870 $Y=435285
X1499 988 1060 263 994 976 1 2 XNR4D2BWP7T $T=305600 451200 1 180 $X=291870 $Y=450965
X1500 992 236 276 1066 1048 1 2 XNR4D2BWP7T $T=296640 459040 0 0 $X=296350 $Y=458805
X1501 1028 1018 285 1069 983 1 2 XNR4D2BWP7T $T=302800 474720 1 0 $X=302510 $Y=470510
X1502 1054 1070 283 1044 1047 1 2 XNR4D2BWP7T $T=319040 443360 0 180 $X=305310 $Y=439150
X1503 1059 1038 289 1072 218 1 2 XNR4D2BWP7T $T=306160 443360 0 0 $X=305870 $Y=443125
X1504 1077 231 287 994 218 1 2 XNR4D2BWP7T $T=321840 451200 1 180 $X=308110 $Y=450965
X1505 92 755 980 1 2 986 MUX2ND1BWP7T $T=229440 474720 1 0 $X=229150 $Y=470510
X1506 771 223 981 1 2 989 MUX2ND1BWP7T $T=232240 435520 1 0 $X=231950 $Y=431310
X1507 92 982 980 1 2 990 MUX2ND1BWP7T $T=232800 451200 0 0 $X=232510 $Y=450965
X1508 975 228 221 1 2 995 MUX2ND1BWP7T $T=233360 459040 1 0 $X=233070 $Y=454830
X1509 1033 908 230 1 2 1037 MUX2ND1BWP7T $T=270880 474720 1 0 $X=270590 $Y=470510
X1510 248 786 1031 1 2 1044 MUX2ND1BWP7T $T=274240 435520 0 0 $X=273950 $Y=435285
X1511 1047 978 260 1 2 1059 MUX2ND1BWP7T $T=296080 435520 1 0 $X=295790 $Y=431310
X1512 1037 986 1040 255 1 2 XNR3D2BWP7T $T=270880 451200 0 0 $X=270590 $Y=450965
X1513 990 1037 1052 267 1 2 XNR3D2BWP7T $T=289920 459040 1 0 $X=289630 $Y=454830
X1514 1045 1047 1062 275 1 2 XNR3D2BWP7T $T=294960 443360 0 0 $X=294670 $Y=443125
X1515 986 1007 1 2 1039 XNR2D1BWP7T $T=268080 451200 1 0 $X=267790 $Y=446990
X1516 958 987 1 2 1041 XNR2D1BWP7T $T=278160 466880 1 180 $X=272830 $Y=466645
X1517 997 1041 1 2 1048 XNR2D1BWP7T $T=277040 474720 1 0 $X=276750 $Y=470510
X1518 262 258 1 2 759 XNR2D1BWP7T $T=294960 419840 1 180 $X=289630 $Y=419605
X1519 252 1045 1 2 1054 XNR2D1BWP7T $T=292160 443360 1 0 $X=291870 $Y=439150
X1520 260 1047 2 1 CKND2BWP7T $T=292720 427680 0 180 $X=290190 $Y=423470
X1521 45 1 2 544 CKND0BWP7T $T=61440 474720 0 180 $X=59470 $Y=470510
X1522 560 1 2 507 CKND0BWP7T $T=62000 435520 1 180 $X=60030 $Y=435285
X1523 29 1 2 686 CKND0BWP7T $T=111280 451200 1 180 $X=109310 $Y=450965
X1524 108 1 2 792 CKND0BWP7T $T=150480 443360 0 0 $X=150190 $Y=443125
X1525 136 1 2 839 CKND0BWP7T $T=174560 419840 0 0 $X=174270 $Y=419605
X1526 150 1 2 797 CKND0BWP7T $T=175120 427680 0 0 $X=174830 $Y=427445
X1527 248 1 2 1031 CKND0BWP7T $T=280400 427680 1 180 $X=278430 $Y=427445
X1528 229 239 1 2 1018 CKXOR2D0BWP7T $T=257440 459040 0 0 $X=257150 $Y=458805
X1529 987 979 1 2 1045 CKXOR2D0BWP7T $T=275360 443360 0 0 $X=275070 $Y=443125
X1530 1033 1041 1 2 1049 CKXOR2D0BWP7T $T=278160 466880 0 0 $X=277870 $Y=466645
X1531 243 229 1007 243 229 2 1 IAO22D1BWP7T $T=262480 443360 1 180 $X=257150 $Y=443125
X1532 223 2 980 969 92 968 1 AOI22D2BWP7T $T=230560 443360 1 180 $X=223550 $Y=443125
X1533 226 2 981 231 771 228 1 AOI22D2BWP7T $T=229440 427680 1 0 $X=229150 $Y=423470
X1534 970 2 980 988 92 216 1 AOI22D2BWP7T $T=229440 459040 0 0 $X=229150 $Y=458805
X1535 229 2 984 994 972 234 1 AOI22D2BWP7T $T=232800 443360 0 0 $X=232510 $Y=443125
X1536 982 2 771 1011 981 723 1 AOI22D2BWP7T $T=249040 459040 0 0 $X=248750 $Y=458805
X1537 241 2 973 1029 1020 1006 1 AOI22D2BWP7T $T=255760 435520 1 0 $X=255470 $Y=431310
X1538 1002 234 229 993 1 2 MUX2ND0BWP7T $T=253520 443360 1 180 $X=248750 $Y=443125
X1539 725 750 706 735 661 2 1 AOI22D0BWP7T $T=133680 451200 1 180 $X=130030 $Y=450965
X1540 891 955 949 960 910 2 1 AOI22D0BWP7T $T=216000 435520 1 0 $X=215710 $Y=431310
X1541 998 991 236 234 229 2 1 AOI22D0BWP7T $T=247920 451200 0 0 $X=247630 $Y=450965
X1542 225 972 230 2 1 992 XNR3D0BWP7T $T=230000 466880 0 0 $X=229710 $Y=466645
X1543 615 1 2 648 CKBD0BWP7T $T=95600 435520 1 180 $X=93070 $Y=435285
X1544 87 1 2 85 CKBD0BWP7T $T=124160 419840 1 180 $X=121630 $Y=419605
X1545 752 1 2 754 CKBD0BWP7T $T=133680 459040 0 0 $X=133390 $Y=458805
X1546 148 1 2 852 CKBD0BWP7T $T=176800 427680 0 0 $X=176510 $Y=427445
X1547 89 1 2 976 CKBD0BWP7T $T=227760 451200 1 0 $X=227470 $Y=446990
X1548 960 833 948 966 2 1 220 AO211D1BWP7T $T=224960 443360 1 0 $X=224670 $Y=439150
X1549 4 2 460 10 1 NR2D1BWP7T $T=21680 443360 1 0 $X=21390 $Y=439150
X1550 17 2 472 16 1 NR2D1BWP7T $T=25600 427680 1 0 $X=25310 $Y=423470
X1551 462 2 487 25 1 NR2D1BWP7T $T=28960 474720 1 0 $X=28670 $Y=470510
X1552 14 2 500 476 1 NR2D1BWP7T $T=44640 466880 0 180 $X=42110 $Y=462670
X1553 545 2 570 459 1 NR2D1BWP7T $T=62000 451200 0 0 $X=61710 $Y=450965
X1554 504 2 576 501 1 NR2D1BWP7T $T=64240 451200 0 0 $X=63950 $Y=450965
X1555 551 2 577 546 1 NR2D1BWP7T $T=64240 459040 1 0 $X=63950 $Y=454830
X1556 461 2 581 33 1 NR2D1BWP7T $T=64800 443360 1 0 $X=64510 $Y=439150
X1557 592 2 598 511 1 NR2D1BWP7T $T=73200 459040 0 180 $X=70670 $Y=454830
X1558 482 2 625 62 1 NR2D1BWP7T $T=87200 419840 1 0 $X=86910 $Y=415630
X1559 60 2 593 573 1 NR2D1BWP7T $T=90000 427680 1 180 $X=87470 $Y=427445
X1560 639 2 597 573 1 NR2D1BWP7T $T=92800 435520 1 180 $X=90270 $Y=435285
X1561 644 2 637 501 1 NR2D1BWP7T $T=93920 451200 0 180 $X=91390 $Y=446990
X1562 45 2 611 638 1 NR2D1BWP7T $T=95600 459040 1 180 $X=93070 $Y=458805
X1563 538 2 658 638 1 NR2D1BWP7T $T=93920 451200 1 0 $X=93630 $Y=446990
X1564 482 2 656 471 1 NR2D1BWP7T $T=96720 466880 1 180 $X=94190 $Y=466645
X1565 73 2 668 71 1 NR2D1BWP7T $T=101760 419840 0 180 $X=99230 $Y=415630
X1566 67 2 673 560 1 NR2D1BWP7T $T=101760 427680 0 0 $X=101470 $Y=427445
X1567 29 2 709 75 1 NR2D1BWP7T $T=111840 443360 1 180 $X=109310 $Y=443125
X1568 3 2 734 731 1 NR2D1BWP7T $T=126960 427680 0 180 $X=124430 $Y=423470
X1569 787 2 776 112 1 NR2D1BWP7T $T=149360 427680 0 0 $X=149070 $Y=427445
X1570 119 2 781 124 1 NR2D1BWP7T $T=153280 443360 0 0 $X=152990 $Y=443125
X1571 127 2 802 768 1 NR2D1BWP7T $T=157200 419840 1 180 $X=154670 $Y=419605
X1572 103 2 788 124 1 NR2D1BWP7T $T=154960 459040 0 0 $X=154670 $Y=458805
X1573 121 2 789 136 1 NR2D1BWP7T $T=164480 427680 1 0 $X=164190 $Y=423470
X1574 827 2 836 125 1 NR2D1BWP7T $T=172880 427680 0 0 $X=172590 $Y=427445
X1575 770 2 862 858 1 NR2D1BWP7T $T=180160 466880 1 0 $X=179870 $Y=462670
X1576 849 2 855 858 1 NR2D1BWP7T $T=185200 466880 0 180 $X=182670 $Y=462670
X1577 857 2 896 181 1 NR2D1BWP7T $T=190240 443360 0 0 $X=189950 $Y=443125
X1578 101 2 892 193 1 NR2D1BWP7T $T=196960 419840 1 0 $X=196670 $Y=415630
X1579 914 2 879 843 1 NR2D1BWP7T $T=199200 435520 0 180 $X=196670 $Y=431310
X1580 195 2 197 892 1 NR2D1BWP7T $T=205920 419840 1 0 $X=205630 $Y=415630
X1581 201 2 853 198 1 NR2D1BWP7T $T=210400 419840 0 180 $X=207870 $Y=415630
X1582 953 2 895 961 1 NR2D1BWP7T $T=218240 459040 0 0 $X=217950 $Y=458805
X1583 964 2 949 954 1 NR2D1BWP7T $T=223840 459040 0 180 $X=221310 $Y=454830
X1584 925 948 896 915 1 2 AOI21D0BWP7T $T=214880 443360 0 0 $X=214590 $Y=443125
X1585 215 959 874 934 1 2 AOI21D0BWP7T $T=219920 427680 1 0 $X=219630 $Y=423470
X1586 484 481 476 9 2 1 474 NR4D1BWP7T $T=30640 451200 1 180 $X=24750 $Y=450965
X1587 486 18 462 9 2 1 14 NR4D1BWP7T $T=30640 466880 1 180 $X=24750 $Y=466645
X1588 499 25 476 490 2 1 20 NR4D1BWP7T $T=43520 443360 1 180 $X=37630 $Y=443125
X1589 523 522 496 29 2 1 18 NR4D1BWP7T $T=50800 451200 1 180 $X=44910 $Y=450965
X1590 527 483 519 513 2 1 460 NR4D1BWP7T $T=51360 435520 1 180 $X=45470 $Y=435285
X1591 532 510 524 459 2 1 505 NR4D1BWP7T $T=52480 459040 0 180 $X=46590 $Y=454830
X1592 561 42 25 541 2 1 545 NR4D1BWP7T $T=59760 443360 1 180 $X=53870 $Y=443125
X1593 557 42 18 548 2 1 509 NR4D1BWP7T $T=61440 443360 0 180 $X=55550 $Y=439150
X1594 558 466 474 509 2 1 40 NR4D1BWP7T $T=62000 435520 0 180 $X=56110 $Y=431310
X1595 565 524 462 542 2 1 555 NR4D1BWP7T $T=63120 459040 1 180 $X=57230 $Y=458805
X1596 571 519 459 553 2 1 547 NR4D1BWP7T $T=64240 459040 0 180 $X=58350 $Y=454830
X1597 567 524 481 554 2 1 511 NR4D1BWP7T $T=64240 466880 0 180 $X=58350 $Y=462670
X1598 587 471 481 555 2 1 14 NR4D1BWP7T $T=68720 466880 1 180 $X=62830 $Y=466645
X1599 564 23 560 574 2 1 490 NR4D1BWP7T $T=69280 427680 1 180 $X=63390 $Y=427445
X1600 584 595 592 566 2 1 522 NR4D1BWP7T $T=72640 474720 0 180 $X=66750 $Y=470510
X1601 640 603 509 621 2 1 629 NR4D1BWP7T $T=91120 466880 0 180 $X=85230 $Y=462670
X1602 650 471 481 63 2 1 516 NR4D1BWP7T $T=94480 466880 1 180 $X=88590 $Y=466645
X1603 664 45 638 513 2 1 639 NR4D1BWP7T $T=97280 435520 0 180 $X=91390 $Y=431310
X1604 652 67 573 606 2 1 73 NR4D1BWP7T $T=94480 427680 0 0 $X=94190 $Y=427445
X1605 665 569 606 663 2 1 636 NR4D1BWP7T $T=101760 443360 0 180 $X=95870 $Y=439150
X1606 662 641 466 75 2 1 14 NR4D1BWP7T $T=97280 435520 0 0 $X=96990 $Y=435285
X1607 649 463 59 638 2 1 690 NR4D1BWP7T $T=101200 435520 1 0 $X=100910 $Y=431310
X1608 769 95 770 763 2 1 93 NR4D1BWP7T $T=144880 427680 1 180 $X=138990 $Y=427445
X1609 772 97 96 91 2 1 94 NR4D1BWP7T $T=146000 419840 0 180 $X=140110 $Y=415630
X1610 765 768 98 777 2 1 793 NR4D1BWP7T $T=142080 435520 0 0 $X=141790 $Y=435285
X1611 803 125 783 793 2 1 114 NR4D1BWP7T $T=157200 435520 0 180 $X=151310 $Y=431310
X1612 801 795 783 794 2 1 805 NR4D1BWP7T $T=151600 466880 1 0 $X=151310 $Y=462670
X1613 813 808 108 816 2 1 146 NR4D1BWP7T $T=163920 466880 1 0 $X=163630 $Y=462670
X1614 821 125 103 823 2 1 146 NR4D1BWP7T $T=165600 459040 0 0 $X=165310 $Y=458805
X1615 829 768 124 824 2 1 835 NR4D1BWP7T $T=168400 466880 0 0 $X=168110 $Y=466645
X1616 779 145 827 814 2 1 155 NR4D1BWP7T $T=168960 427680 1 0 $X=168670 $Y=423470
X1617 840 125 827 151 2 1 820 NR4D1BWP7T $T=176240 466880 0 180 $X=170350 $Y=462670
X1618 844 843 145 834 2 1 811 NR4D1BWP7T $T=178480 443360 0 180 $X=172590 $Y=439150
X1619 846 143 809 812 2 1 838 NR4D1BWP7T $T=179040 451200 1 180 $X=173150 $Y=450965
X1620 845 124 143 849 2 1 800 NR4D1BWP7T $T=174000 466880 0 0 $X=173710 $Y=466645
X1621 874 171 860 143 2 1 121 NR4D1BWP7T $T=186880 427680 0 180 $X=180990 $Y=423470
X1622 886 876 809 856 2 1 820 NR4D1BWP7T $T=188560 443360 1 180 $X=182670 $Y=443125
X1623 890 883 808 869 2 1 820 NR4D1BWP7T $T=190240 459040 0 180 $X=184350 $Y=454830
X1624 901 184 897 868 2 1 861 NR4D1BWP7T $T=194160 451200 1 180 $X=188270 $Y=450965
X1625 847 182 145 906 2 1 178 NR4D1BWP7T $T=190240 427680 1 0 $X=189950 $Y=423470
X1626 907 169 900 865 2 1 902 NR4D1BWP7T $T=191360 435520 0 0 $X=191070 $Y=435285
X1627 894 843 187 870 2 1 181 NR4D1BWP7T $T=196960 459040 1 180 $X=191070 $Y=458805
X1628 918 182 145 906 2 1 178 NR4D1BWP7T $T=199200 427680 1 180 $X=193310 $Y=427445
X1629 938 170 208 201 2 1 98 NR4D1BWP7T $T=216000 419840 0 180 $X=210110 $Y=415630
X1630 944 176 201 854 2 1 210 NR4D1BWP7T $T=224400 419840 0 180 $X=218510 $Y=415630
X1631 957 916 956 2 1 963 AN3D1BWP7T $T=218240 443360 1 0 $X=217950 $Y=439150
X1632 880 2 871 840 855 801 1 AOI31D2BWP7T $T=188000 466880 1 180 $X=180990 $Y=466645
X1633 880 2 889 185 882 846 1 AOI31D2BWP7T $T=195840 466880 1 180 $X=188830 $Y=466645
X1634 915 2 873 796 766 192 1 AOI31D2BWP7T $T=199200 459040 0 180 $X=192190 $Y=454830
X1635 884 2 899 191 894 898 1 AOI31D2BWP7T $T=199200 466880 0 180 $X=192190 $Y=462670
X1636 934 2 913 927 922 829 1 AOI31D2BWP7T $T=212640 466880 1 180 $X=205630 $Y=466645
X1637 934 2 937 875 796 901 1 AOI31D2BWP7T $T=214320 466880 0 180 $X=207310 $Y=462670
X1638 884 2 950 927 194 935 1 AOI31D2BWP7T $T=217680 474720 0 180 $X=210670 $Y=470510
X1639 915 2 962 918 928 213 1 AOI31D2BWP7T $T=224960 435520 1 180 $X=217950 $Y=435285
X1640 939 921 959 940 2 1 965 OR4D1BWP7T $T=217680 443360 0 0 $X=217390 $Y=443125
X1641 642 671 578 608 1 2 694 OA31D0BWP7T $T=103440 466880 0 0 $X=103150 $Y=466645
X1642 712 485 635 735 1 2 737 OA31D0BWP7T $T=122480 466880 0 0 $X=122190 $Y=466645
X1643 691 88 485 706 1 2 739 OA31D0BWP7T $T=123600 459040 0 0 $X=123310 $Y=458805
X1644 546 516 749 677 1 2 753 OA31D0BWP7T $T=131440 466880 1 0 $X=131150 $Y=462670
X1645 135 212 214 960 1 2 945 OA31D0BWP7T $T=217680 419840 0 0 $X=217390 $Y=419605
X1646 17 2 459 3 4 1 AOI21D2BWP7T $T=26160 459040 0 180 $X=20830 $Y=454830
X1647 524 2 550 31 464 1 AOI21D2BWP7T $T=59200 466880 1 180 $X=53870 $Y=466645
X1648 947 2 958 951 949 1 AOI21D2BWP7T $T=216560 451200 0 0 $X=216270 $Y=450965
X1649 24 1 473 19 2 ND2D1BWP7T $T=31200 435520 0 180 $X=28670 $Y=431310
X1650 488 1 493 464 2 ND2D1BWP7T $T=39040 427680 0 0 $X=38750 $Y=427445
X1651 7 1 494 495 2 ND2D1BWP7T $T=40160 419840 0 0 $X=39870 $Y=419605
X1652 488 1 497 480 2 ND2D1BWP7T $T=40720 435520 1 0 $X=40430 $Y=431310
X1653 488 1 503 495 2 ND2D1BWP7T $T=42400 419840 0 0 $X=42110 $Y=419605
X1654 495 1 492 27 2 ND2D1BWP7T $T=42960 419840 1 0 $X=42670 $Y=415630
X1655 32 1 22 27 2 ND2D1BWP7T $T=49680 419840 0 180 $X=47150 $Y=415630
X1656 32 1 517 7 2 ND2D1BWP7T $T=49680 419840 1 180 $X=47150 $Y=419605
X1657 38 1 34 480 2 ND2D1BWP7T $T=53040 427680 0 180 $X=50510 $Y=423470
X1658 495 1 35 31 2 ND2D1BWP7T $T=53600 419840 0 180 $X=51070 $Y=415630
X1659 38 1 531 495 2 ND2D1BWP7T $T=55840 427680 0 180 $X=53310 $Y=423470
X1660 26 1 40 493 2 ND2D1BWP7T $T=56960 419840 0 180 $X=54430 $Y=415630
X1661 43 1 548 502 2 ND2D1BWP7T $T=59200 427680 0 180 $X=56670 $Y=423470
X1662 41 1 521 480 2 ND2D1BWP7T $T=57520 419840 0 0 $X=57230 $Y=419605
X1663 517 1 547 44 2 ND2D1BWP7T $T=58640 451200 1 0 $X=58350 $Y=446990
X1664 38 1 549 464 2 ND2D1BWP7T $T=59200 427680 0 0 $X=58910 $Y=427445
X1665 41 1 556 495 2 ND2D1BWP7T $T=59760 419840 0 0 $X=59470 $Y=419605
X1666 495 1 559 19 2 ND2D1BWP7T $T=60320 427680 1 0 $X=60030 $Y=423470
X1667 19 1 26 49 2 ND2D1BWP7T $T=61440 419840 1 0 $X=61150 $Y=415630
X1668 556 1 563 527 2 ND2D1BWP7T $T=63680 443360 0 180 $X=61150 $Y=439150
X1669 544 1 566 44 2 ND2D1BWP7T $T=61440 474720 1 0 $X=61150 $Y=470510
X1670 47 1 518 495 2 ND2D1BWP7T $T=64800 419840 1 180 $X=62270 $Y=419605
X1671 494 1 555 575 2 ND2D1BWP7T $T=63120 459040 0 0 $X=62830 $Y=458805
X1672 24 1 572 7 2 ND2D1BWP7T $T=68720 419840 0 180 $X=66190 $Y=415630
X1673 7 1 575 49 2 ND2D1BWP7T $T=70960 419840 0 180 $X=68430 $Y=415630
X1674 47 1 591 480 2 ND2D1BWP7T $T=68720 419840 0 0 $X=68430 $Y=419605
X1675 571 1 599 550 2 ND2D1BWP7T $T=70400 459040 0 0 $X=70110 $Y=458805
X1676 38 1 582 49 2 ND2D1BWP7T $T=73200 419840 1 180 $X=70670 $Y=419605
X1677 601 1 528 521 2 ND2D1BWP7T $T=73200 443360 0 180 $X=70670 $Y=439150
X1678 575 1 53 48 2 ND2D1BWP7T $T=79920 419840 1 0 $X=79630 $Y=415630
X1679 34 1 614 625 2 ND2D1BWP7T $T=83280 443360 0 0 $X=82990 $Y=443125
X1680 497 1 594 593 2 ND2D1BWP7T $T=83840 435520 0 0 $X=83550 $Y=435285
X1681 492 1 509 630 2 ND2D1BWP7T $T=86080 466880 0 0 $X=85790 $Y=466645
X1682 22 1 636 26 2 ND2D1BWP7T $T=88880 419840 0 0 $X=88590 $Y=419605
X1683 559 1 681 68 2 ND2D1BWP7T $T=105120 435520 1 180 $X=102590 $Y=435285
X1684 7 1 633 464 2 ND2D1BWP7T $T=107360 427680 0 180 $X=104830 $Y=423470
X1685 580 1 730 596 2 ND2D1BWP7T $T=126400 443360 0 180 $X=123870 $Y=439150
X1686 757 1 744 762 2 ND2D1BWP7T $T=138160 451200 1 0 $X=137870 $Y=446990
X1687 782 1 91 789 2 ND2D1BWP7T $T=147680 451200 1 0 $X=147390 $Y=446990
X1688 113 1 774 118 2 ND2D1BWP7T $T=151040 451200 1 0 $X=150750 $Y=446990
X1689 115 1 114 120 2 ND2D1BWP7T $T=156080 427680 1 180 $X=153550 $Y=427445
X1690 122 1 793 130 2 ND2D1BWP7T $T=154400 443360 1 0 $X=154110 $Y=439150
X1691 131 1 807 123 2 ND2D1BWP7T $T=163920 419840 0 0 $X=163630 $Y=419605
X1692 129 1 806 784 2 ND2D1BWP7T $T=163920 451200 0 0 $X=163630 $Y=450965
X1693 134 1 814 137 2 ND2D1BWP7T $T=166720 427680 1 0 $X=166430 $Y=423470
X1694 819 1 135 781 2 ND2D1BWP7T $T=169520 443360 0 180 $X=166990 $Y=439150
X1695 128 1 820 142 2 ND2D1BWP7T $T=167840 443360 0 0 $X=167550 $Y=443125
X1696 161 1 848 803 2 ND2D1BWP7T $T=179600 435520 0 180 $X=177070 $Y=431310
X1697 139 1 861 132 2 ND2D1BWP7T $T=180160 419840 0 0 $X=179870 $Y=419605
X1698 867 1 858 141 2 ND2D1BWP7T $T=182960 443360 1 180 $X=180430 $Y=443125
X1699 175 1 865 852 2 ND2D1BWP7T $T=184080 427680 1 180 $X=181550 $Y=427445
X1700 168 1 831 144 2 ND2D1BWP7T $T=184640 451200 1 180 $X=182110 $Y=450965
X1701 792 1 902 904 2 ND2D1BWP7T $T=192480 443360 1 0 $X=192190 $Y=439150
X1702 839 1 885 186 2 ND2D1BWP7T $T=195840 419840 1 180 $X=193310 $Y=419605
X1703 917 1 906 137 2 ND2D1BWP7T $T=198080 427680 0 180 $X=195550 $Y=423470
X1704 194 1 900 828 2 ND2D1BWP7T $T=199200 435520 1 180 $X=196670 $Y=435285
X1705 953 1 934 954 2 ND2D1BWP7T $T=216000 459040 0 0 $X=215710 $Y=458805
X1706 473 1 468 13 2 470 8 OAI211D1BWP7T $T=26720 466880 0 180 $X=23070 $Y=462670
X1707 670 1 617 640 2 683 687 OAI211D1BWP7T $T=102320 466880 1 0 $X=102030 $Y=462670
X1708 61 1 56 708 2 700 82 OAI211D1BWP7T $T=108480 427680 0 0 $X=108190 $Y=427445
X1709 686 1 668 722 2 663 13 OAI211D1BWP7T $T=111840 435520 0 0 $X=111550 $Y=435285
X1710 526 1 709 708 2 725 13 OAI211D1BWP7T $T=111840 443360 0 0 $X=111550 $Y=443125
X1711 668 1 580 728 2 721 3 OAI211D1BWP7T $T=121920 435520 0 0 $X=121630 $Y=435285
X1712 515 1 596 83 2 732 10 OAI211D1BWP7T $T=122480 427680 0 0 $X=122190 $Y=427445
X1713 779 1 776 101 2 763 99 OAI211D1BWP7T $T=147680 419840 1 180 $X=144030 $Y=419605
X1714 149 1 152 154 2 825 156 OAI211D1BWP7T $T=171200 419840 0 0 $X=170910 $Y=419605
X1715 797 1 161 163 2 856 156 OAI211D1BWP7T $T=176240 427680 1 0 $X=175950 $Y=423470
X1716 839 1 919 101 2 914 156 OAI211D1BWP7T $T=205920 427680 1 0 $X=205630 $Y=423470
X1717 888 1 943 821 2 947 934 OAI211D1BWP7T $T=212640 459040 0 0 $X=212350 $Y=458805
X1718 924 1 955 211 2 971 884 OAI211D1BWP7T $T=216000 427680 0 0 $X=215710 $Y=427445
X1719 25 2 510 483 471 1 515 NR4D2BWP7T $T=50800 466880 1 180 $X=37630 $Y=466645
X1720 491 2 469 520 483 1 526 NR4D2BWP7T $T=40160 459040 0 0 $X=39870 $Y=458805
X1721 607 2 55 595 553 1 646 NR4D2BWP7T $T=79920 474720 1 0 $X=79630 $Y=470510
X1722 811 2 807 121 876 1 875 NR4D2BWP7T $T=175120 435520 0 0 $X=174830 $Y=435285
X1723 950 2 871 962 937 1 979 NR4D2BWP7T $T=228320 466880 1 180 $X=215150 $Y=466645
X1724 165 2 838 826 1 NR2XD0BWP7T $T=180720 443360 0 180 $X=178190 $Y=439150
X1725 953 2 954 936 1 NR2XD0BWP7T $T=217680 459040 0 180 $X=215150 $Y=454830
X1726 880 778 872 884 2 1 929 OA22D0BWP7T $T=205920 443360 1 0 $X=205630 $Y=439150
X1727 884 946 830 915 2 1 956 OA22D0BWP7T $T=213760 435520 0 0 $X=213470 $Y=435285
X1728 508 1 30 34 531 538 2 ND4D1BWP7T $T=50800 451200 0 0 $X=50510 $Y=450965
X1729 518 1 493 37 517 542 2 ND4D1BWP7T $T=51360 419840 0 0 $X=51070 $Y=419605
X1730 34 1 537 500 502 552 2 ND4D1BWP7T $T=52480 451200 1 0 $X=52190 $Y=446990
X1731 588 1 503 584 468 583 2 ND4D1BWP7T $T=69840 459040 1 180 $X=65630 $Y=458805
X1732 497 1 52 589 54 615 2 ND4D1BWP7T $T=79920 435520 0 0 $X=79630 $Y=435285
X1733 565 1 611 609 596 607 2 ND4D1BWP7T $T=79920 459040 0 0 $X=79630 $Y=458805
X1734 582 1 588 589 492 628 2 ND4D1BWP7T $T=80480 451200 0 0 $X=80190 $Y=450965
X1735 591 1 48 576 58 627 2 ND4D1BWP7T $T=82720 435520 1 0 $X=82430 $Y=431310
X1736 559 1 631 58 581 629 2 ND4D1BWP7T $T=90000 435520 1 180 $X=85790 $Y=435285
X1737 508 1 662 656 550 671 2 ND4D1BWP7T $T=96720 466880 0 0 $X=96430 $Y=466645
X1738 113 1 117 116 106 791 2 ND4D1BWP7T $T=154400 419840 0 180 $X=150190 $Y=415630
X1739 129 1 115 789 111 800 2 ND4D1BWP7T $T=157200 451200 1 180 $X=152990 $Y=450965
X1740 804 1 129 784 141 811 2 ND4D1BWP7T $T=164480 451200 1 0 $X=164190 $Y=446990
X1741 139 1 115 122 132 812 2 ND4D1BWP7T $T=166160 419840 0 0 $X=165870 $Y=419605
X1742 772 1 822 826 819 833 2 ND4D1BWP7T $T=168960 435520 0 0 $X=168670 $Y=435285
X1743 128 1 117 828 152 816 2 ND4D1BWP7T $T=170080 443360 0 0 $X=169790 $Y=443125
X1744 159 1 149 158 802 834 2 ND4D1BWP7T $T=177920 419840 0 180 $X=173710 $Y=415630
X1745 128 1 160 847 851 854 2 ND4D1BWP7T $T=176240 419840 0 0 $X=175950 $Y=419605
X1746 209 1 197 196 927 951 2 ND4D1BWP7T $T=213760 419840 0 0 $X=213470 $Y=419605
X1747 520 594 670 674 677 1 2 OAI31D1BWP7T $T=98400 466880 1 0 $X=98110 $Y=462670
X1748 606 470 684 685 608 1 2 OAI31D1BWP7T $T=102880 451200 0 0 $X=102590 $Y=450965
X1749 624 698 696 643 677 1 2 OAI31D1BWP7T $T=109600 459040 0 180 $X=105390 $Y=454830
X1750 700 671 697 583 677 1 2 OAI31D1BWP7T $T=109600 466880 0 180 $X=105390 $Y=462670
X1751 698 603 711 692 608 1 2 OAI31D1BWP7T $T=109600 459040 1 0 $X=109310 $Y=454830
X1752 657 678 720 603 706 1 2 OAI31D1BWP7T $T=111280 451200 0 0 $X=110990 $Y=450965
X1753 553 712 719 669 706 1 2 OAI31D1BWP7T $T=115200 466880 0 180 $X=110990 $Y=462670
X1754 553 563 727 714 706 1 2 OAI31D1BWP7T $T=125840 451200 1 180 $X=121630 $Y=450965
X1755 730 672 729 530 735 1 2 OAI31D1BWP7T $T=124160 451200 1 0 $X=123870 $Y=446990
X1756 628 546 752 675 608 1 2 OAI31D1BWP7T $T=131440 459040 1 0 $X=131150 $Y=454830
X1757 808 858 888 791 895 1 2 OAI31D1BWP7T $T=187440 459040 0 0 $X=187150 $Y=458805
X1758 112 199 924 923 936 1 2 OAI31D1BWP7T $T=207600 427680 0 0 $X=207310 $Y=427445
X1759 206 848 943 942 936 1 2 OAI31D1BWP7T $T=212080 427680 0 0 $X=211790 $Y=427445
X1760 699 543 741 745 746 1 2 AOI31D0BWP7T $T=128640 443360 1 0 $X=128350 $Y=439150
X1761 200 890 785 926 915 1 2 AOI31D0BWP7T $T=209840 459040 0 180 $X=206190 $Y=454830
X1762 844 930 205 933 880 1 2 AOI31D0BWP7T $T=209280 443360 0 0 $X=208990 $Y=443125
X1763 203 194 928 939 884 1 2 AOI31D0BWP7T $T=210400 435520 0 0 $X=210110 $Y=435285
X1764 905 194 886 940 915 1 2 AOI31D0BWP7T $T=211520 451200 1 0 $X=211230 $Y=446990
X1765 633 1 26 68 2 667 ND3D0BWP7T $T=95600 419840 0 0 $X=95310 $Y=419605
X1766 634 1 69 658 2 672 ND3D0BWP7T $T=96160 451200 1 0 $X=95870 $Y=446990
X1767 917 1 938 890 2 206 ND3D0BWP7T $T=210960 427680 1 0 $X=210670 $Y=423470
X1768 9 1 2 20 472 478 23 NR4D0BWP7T $T=27840 427680 1 0 $X=27550 $Y=423470
X1769 460 1 2 33 11 533 519 NR4D0BWP7T $T=49680 443360 1 0 $X=49390 $Y=439150
X1770 525 1 2 511 11 535 463 NR4D0BWP7T $T=53040 459040 0 0 $X=52750 $Y=458805
X1771 45 1 2 9 14 562 471 NR4D0BWP7T $T=63120 466880 1 180 $X=59470 $Y=466645
X1772 614 1 2 599 481 613 462 NR4D0BWP7T $T=83280 466880 0 180 $X=79630 $Y=462670
X1773 627 1 2 623 509 622 603 NR4D0BWP7T $T=87200 443360 0 180 $X=83550 $Y=439150
X1774 636 1 2 639 505 634 610 NR4D0BWP7T $T=92240 443360 0 180 $X=88590 $Y=439150
X1775 648 1 2 599 462 645 638 NR4D0BWP7T $T=93360 459040 1 180 $X=89710 $Y=458805
X1776 552 1 2 678 516 699 681 NR4D0BWP7T $T=106240 443360 1 0 $X=105950 $Y=439150
X1777 612 1 2 672 586 705 690 NR4D0BWP7T $T=107360 451200 1 0 $X=107070 $Y=446990
X1778 721 1 2 678 638 717 463 NR4D0BWP7T $T=112960 443360 0 180 $X=109310 $Y=439150
X1779 666 1 2 485 534 733 546 NR4D0BWP7T $T=122480 474720 1 0 $X=122190 $Y=470510
X1780 627 1 2 734 14 736 690 NR4D0BWP7T $T=126960 435520 0 180 $X=123310 $Y=431310
X1781 726 1 2 590 563 740 14 NR4D0BWP7T $T=126960 451200 0 0 $X=126670 $Y=450965
X1782 800 1 2 838 831 842 820 NR4D0BWP7T $T=177360 459040 0 180 $X=173710 $Y=454830
X1783 167 1 2 807 820 866 848 NR4D0BWP7T $T=184080 443360 0 180 $X=180430 $Y=439150
X1784 180 1 2 173 176 878 169 NR4D0BWP7T $T=190240 419840 0 180 $X=186590 $Y=415630
X1785 885 1 2 865 835 893 790 NR4D0BWP7T $T=191360 435520 1 180 $X=187710 $Y=435285
X1786 805 1 2 902 155 905 188 NR4D0BWP7T $T=191920 451200 1 0 $X=191630 $Y=446990
X1787 202 1 2 188 809 925 897 NR4D0BWP7T $T=210400 451200 0 180 $X=206750 $Y=446990
X1788 926 1 2 877 933 932 945 NR4D0BWP7T $T=209840 459040 1 0 $X=209550 $Y=454830
X1789 6 11 2 465 1 NR2D2BWP7T $T=30640 443360 0 180 $X=26430 $Y=439150
X1790 472 474 2 498 1 NR2D2BWP7T $T=39040 427680 1 0 $X=38750 $Y=423470
X1791 461 569 2 580 1 NR2D2BWP7T $T=65360 443360 0 0 $X=65070 $Y=443125
X1792 81 10 2 560 1 NR2D2BWP7T $T=111280 419840 1 180 $X=107070 $Y=419605
X1793 859 920 2 927 1 NR2D2BWP7T $T=208160 419840 0 0 $X=207870 $Y=419605
X1794 580 572 503 521 2 1 604 AN4D1BWP7T $T=67600 435520 0 0 $X=67310 $Y=435285
X1795 487 581 649 508 2 1 655 AN4D1BWP7T $T=91680 466880 1 0 $X=91390 $Y=462670
X1796 713 719 711 697 2 1 723 AN4D1BWP7T $T=111280 459040 0 0 $X=110990 $Y=458805
X1797 727 729 696 684 2 1 89 AN4D1BWP7T $T=123040 459040 1 0 $X=122750 $Y=454830
X1798 132 142 815 140 2 1 822 AN4D1BWP7T $T=166720 427680 0 0 $X=166430 $Y=427445
X1799 118 126 157 867 2 1 887 AN4D1BWP7T $T=183520 451200 1 0 $X=183230 $Y=446990
X1800 111 875 919 134 2 1 928 AN4D1BWP7T $T=206480 435520 0 0 $X=206190 $Y=435285
X1801 564 1 2 568 BUFFD0BWP7T $T=61440 427680 0 0 $X=61150 $Y=427445
X1802 567 1 2 579 BUFFD0BWP7T $T=64240 466880 1 0 $X=63950 $Y=462670
X1803 613 1 2 620 BUFFD0BWP7T $T=83280 466880 1 0 $X=82990 $Y=462670
X1804 765 1 2 766 BUFFD0BWP7T $T=141520 435520 1 0 $X=141230 $Y=431310
X1805 866 1 2 872 BUFFD0BWP7T $T=184080 443360 1 0 $X=183790 $Y=439150
X1806 785 1 2 922 BUFFD0BWP7T $T=205920 474720 1 0 $X=205630 $Y=470510
X1807 717 695 710 489 687 2 1 AOI31D1BWP7T $T=114640 451200 0 180 $X=110430 $Y=446990
X1808 568 682 738 689 746 2 1 AOI31D1BWP7T $T=127520 443360 0 0 $X=127230 $Y=443125
X1809 813 862 877 882 884 2 1 AOI31D1BWP7T $T=185200 466880 1 0 $X=184910 $Y=462670
X1810 845 196 921 191 880 2 1 AOI31D1BWP7T $T=205920 459040 0 0 $X=205630 $Y=458805
X1811 30 1 518 521 493 525 2 ND4D0BWP7T $T=47440 427680 1 0 $X=47150 $Y=423470
X1812 529 1 507 503 465 541 2 ND4D0BWP7T $T=53040 435520 0 0 $X=52750 $Y=435285
X1813 549 1 46 507 517 554 2 ND4D0BWP7T $T=64240 451200 0 180 $X=60590 $Y=446990
X1814 559 1 503 572 536 574 2 ND4D0BWP7T $T=62000 435520 0 0 $X=61710 $Y=435285
X1815 575 1 556 561 597 605 2 ND4D0BWP7T $T=69280 443360 0 0 $X=68990 $Y=443125
X1816 556 1 52 609 598 612 2 ND4D0BWP7T $T=79920 443360 0 0 $X=79630 $Y=443125
X1817 22 1 591 57 43 626 2 ND4D0BWP7T $T=82160 419840 1 0 $X=81870 $Y=415630
X1818 22 1 588 54 43 619 2 ND4D0BWP7T $T=82160 419840 0 0 $X=81870 $Y=419605
X1819 540 1 51 616 56 621 2 ND4D0BWP7T $T=82160 466880 0 0 $X=81870 $Y=466645
X1820 601 1 622 625 632 647 2 ND4D0BWP7T $T=86640 443360 0 0 $X=86350 $Y=443125
X1821 587 1 61 536 616 635 2 ND4D0BWP7T $T=86640 459040 1 0 $X=86350 $Y=454830
X1822 591 1 46 637 598 642 2 ND4D0BWP7T $T=88320 451200 1 0 $X=88030 $Y=446990
X1823 65 1 499 64 616 657 2 ND4D0BWP7T $T=95600 443360 0 180 $X=91950 $Y=439150
X1824 604 1 600 654 658 661 2 ND4D0BWP7T $T=93920 451200 0 0 $X=93630 $Y=450965
X1825 653 1 665 69 550 675 2 ND4D0BWP7T $T=96720 459040 1 0 $X=96430 $Y=454830
X1826 484 1 70 665 637 669 2 ND4D0BWP7T $T=97280 451200 0 0 $X=96990 $Y=450965
X1827 72 1 654 577 673 676 2 ND4D0BWP7T $T=98400 459040 0 0 $X=98110 $Y=458805
X1828 601 1 591 680 597 691 2 ND4D0BWP7T $T=101200 451200 1 0 $X=100910 $Y=446990
X1829 72 1 620 465 680 688 2 ND4D0BWP7T $T=101760 459040 0 0 $X=101470 $Y=458805
X1830 686 1 645 577 536 679 2 ND4D0BWP7T $T=105680 459040 0 180 $X=102030 $Y=454830
X1831 633 1 467 77 61 692 2 ND4D0BWP7T $T=104000 419840 0 0 $X=103710 $Y=419605
X1832 579 1 558 695 651 701 2 ND4D0BWP7T $T=106240 443360 0 0 $X=105950 $Y=443125
X1833 559 1 631 707 79 714 2 ND4D0BWP7T $T=108480 435520 0 0 $X=108190 $Y=435285
X1834 682 1 580 709 557 726 2 ND4D0BWP7T $T=125840 443360 1 180 $X=122190 $Y=443125
X1835 782 1 105 788 111 794 2 ND4D0BWP7T $T=148240 459040 0 0 $X=147950 $Y=458805
X1836 797 1 792 782 115 787 2 ND4D0BWP7T $T=154400 443360 0 180 $X=150750 $Y=439150
X1837 131 1 134 784 137 799 2 ND4D0BWP7T $T=163920 435520 0 0 $X=163630 $Y=435285
X1838 133 1 784 798 140 817 2 ND4D0BWP7T $T=164480 435520 1 0 $X=164190 $Y=431310
X1839 128 1 120 144 153 824 2 ND4D0BWP7T $T=170080 451200 0 0 $X=169790 $Y=450965
X1840 120 1 842 852 853 823 2 ND4D0BWP7T $T=176800 459040 0 0 $X=176510 $Y=458805
X1841 157 1 164 788 855 857 2 ND4D0BWP7T $T=177360 451200 1 0 $X=177070 $Y=446990
X1842 115 1 138 144 828 868 2 ND4D0BWP7T $T=181280 459040 1 0 $X=180990 $Y=454830
X1843 138 1 126 144 853 870 2 ND4D0BWP7T $T=182400 459040 0 0 $X=182110 $Y=458805
X1844 174 1 878 166 853 891 2 ND4D0BWP7T $T=186880 427680 1 0 $X=186590 $Y=423470
X1845 168 1 903 190 766 910 2 ND4D0BWP7T $T=193600 435520 1 0 $X=193310 $Y=431310
X1846 887 1 886 851 196 923 2 ND4D0BWP7T $T=205920 443360 0 0 $X=205630 $Y=443125
X1847 482 1 492 2 475 491 IND3D1BWP7T $T=41280 435520 1 180 $X=37630 $Y=435285
X1848 155 1 815 2 168 183 IND3D1BWP7T $T=190240 419840 1 0 $X=189950 $Y=415630
X1849 165 1 153 2 134 897 IND3D1BWP7T $T=195280 451200 1 0 $X=194990 $Y=446990
X1850 732 600 627 2 1 NR2D1P5BWP7T $T=129200 435520 1 180 $X=124990 $Y=435285
X1851 84 758 80 2 1 NR2D1P5BWP7T $T=137600 419840 0 0 $X=137310 $Y=419605
X1852 892 815 860 2 1 NR2D1P5BWP7T $T=191360 427680 1 180 $X=187150 $Y=427445
X1853 883 828 187 2 1 NR2D1P5BWP7T $T=194160 451200 0 0 $X=193870 $Y=450965
X1854 99 189 134 2 1 904 OA21D0BWP7T $T=196960 419840 0 180 $X=193310 $Y=415630
X1855 536 2 45 14 60 653 1 INR4D0BWP7T $T=96720 459040 0 180 $X=91950 $Y=454830
X1856 879 2 114 181 900 903 1 INR4D0BWP7T $T=189120 435520 1 0 $X=188830 $Y=431310
X1857 815 2 827 178 177 911 1 INR4D0BWP7T $T=192480 443360 0 0 $X=192190 $Y=443125
X1858 155 1 815 168 2 849 IND3D0BWP7T $T=191920 451200 0 180 $X=188270 $Y=446990
X1859 476 1 504 29 468 2 NR3D1BWP7T $T=45200 459040 0 180 $X=40430 $Y=454830
X1860 644 1 53 626 651 2 NR3D1BWP7T $T=90000 419840 1 0 $X=89710 $Y=415630
X1861 74 1 615 667 682 2 NR3D1BWP7T $T=98400 419840 0 0 $X=98110 $Y=419605
X1862 482 1 534 730 689 2 NR3D1BWP7T $T=125280 466880 1 0 $X=124990 $Y=462670
X1863 91 1 774 775 785 2 NR3D1BWP7T $T=144880 451200 0 0 $X=144590 $Y=450965
X1864 860 1 831 179 882 2 NR3D1BWP7T $T=192480 443360 0 180 $X=187710 $Y=439150
X1865 9 1 584 600 602 517 2 IND4D0BWP7T $T=69280 466880 0 0 $X=68990 $Y=466645
X1866 522 1 536 576 624 601 2 IND4D0BWP7T $T=82720 459040 1 0 $X=82430 $Y=454830
X1867 60 1 570 632 643 582 2 IND4D0BWP7T $T=87200 451200 0 0 $X=86910 $Y=450965
X1868 681 1 651 54 674 65 2 IND4D0BWP7T $T=105680 443360 0 180 $X=101470 $Y=439150
X1869 76 1 597 651 685 689 2 IND4D0BWP7T $T=102320 443360 0 0 $X=102030 $Y=443125
X1870 103 1 106 784 777 110 2 IND4D0BWP7T $T=146560 427680 1 0 $X=146270 $Y=423470
X1871 812 1 815 804 818 113 2 IND4D0BWP7T $T=170080 451200 1 180 $X=165870 $Y=450965
X1872 176 1 126 157 869 867 2 IND4D0BWP7T $T=188560 451200 1 180 $X=184350 $Y=450965
X1873 177 1 879 117 881 784 2 IND4D0BWP7T $T=189120 435520 0 180 $X=184910 $Y=431310
X1874 509 1 500 514 530 517 2 IND4D1BWP7T $T=44640 451200 1 0 $X=44350 $Y=446990
X1875 11 1 35 549 551 494 2 IND4D1BWP7T $T=54160 459040 1 0 $X=53870 $Y=454830
X1876 594 1 571 35 578 575 2 IND4D1BWP7T $T=70960 459040 0 180 $X=66190 $Y=454830
X1877 592 1 652 630 666 68 2 IND4D1BWP7T $T=94480 474720 1 0 $X=94190 $Y=470510
X1878 143 1 138 782 810 133 2 IND4D1BWP7T $T=168400 466880 1 180 $X=163630 $Y=466645
X1879 858 1 162 828 838 802 2 IND4D1BWP7T $T=179600 443360 1 180 $X=174830 $Y=443125
X1880 170 1 132 141 859 117 2 IND4D1BWP7T $T=184640 419840 0 180 $X=179870 $Y=415630
X1881 885 1 836 172 173 126 2 IND4D1BWP7T $T=188560 419840 1 180 $X=183790 $Y=419605
X1882 873 2 889 899 913 1 908 NR4D3BWP7T $T=183520 474720 1 0 $X=183230 $Y=470510
X1883 647 648 644 569 2 1 660 OR4D0BWP7T $T=92800 443360 0 0 $X=92510 $Y=443125
X1884 818 806 150 827 2 1 832 OR4D0BWP7T $T=169520 459040 1 0 $X=169230 $Y=454830
X1885 9 6 469 467 26 1 2 INR4D1BWP7T $T=22240 419840 0 0 $X=21950 $Y=419605
X1886 496 501 20 477 473 1 2 INR4D1BWP7T $T=45200 451200 1 180 $X=38190 $Y=450965
X1887 95 795 121 798 128 1 2 INR4D1BWP7T $T=150480 427680 1 0 $X=150190 $Y=423470
X1888 825 790 817 830 826 1 2 INR4D1BWP7T $T=169520 435520 1 0 $X=169230 $Y=431310
X1889 113 807 1 147 148 2 INR3D1BWP7T $T=166720 419840 1 0 $X=166430 $Y=415630
X1890 122 108 111 2 1 INR2D2BWP7T $T=153840 459040 0 180 $X=149070 $Y=454830
X1891 458 2 461 1 13 NR2XD1BWP7T $T=21120 451200 0 0 $X=20830 $Y=450965
X1892 458 2 462 1 3 NR2XD1BWP7T $T=21120 466880 0 0 $X=20830 $Y=466645
X1893 8 2 463 1 16 NR2XD1BWP7T $T=21680 427680 1 0 $X=21390 $Y=423470
X1894 3 2 466 1 10 NR2XD1BWP7T $T=22800 435520 0 0 $X=22510 $Y=435285
X1895 12 2 6 1 16 NR2XD1BWP7T $T=23920 427680 0 0 $X=23630 $Y=427445
X1896 21 2 474 1 10 NR2XD1BWP7T $T=42400 419840 0 180 $X=38190 $Y=415630
X1897 42 2 596 1 463 NR2XD1BWP7T $T=69280 427680 0 0 $X=68990 $Y=427445
X1898 10 2 644 1 13 NR2XD1BWP7T $T=98960 419840 0 180 $X=94750 $Y=415630
X1899 728 2 90 1 742 NR2XD1BWP7T $T=134800 419840 0 180 $X=130590 $Y=415630
X1900 759 2 706 1 757 NR2XD1BWP7T $T=142080 443360 0 180 $X=137870 $Y=439150
X1901 757 2 608 1 762 NR2XD1BWP7T $T=144320 451200 0 180 $X=140110 $Y=446990
X1902 101 2 783 1 109 NR2XD1BWP7T $T=146560 419840 1 0 $X=146270 $Y=415630
X1903 12 1 475 19 2 IND2D1BWP7T $T=26160 435520 1 0 $X=25870 $Y=431310
X1904 481 1 522 30 2 IND2D1BWP7T $T=49680 466880 1 0 $X=49390 $Y=462670
X1905 547 1 545 39 2 IND2D1BWP7T $T=57520 451200 1 180 $X=54430 $Y=450965
X1906 774 1 104 781 2 IND2D1BWP7T $T=145440 443360 0 0 $X=145150 $Y=443125
X1907 737 694 739 753 2 1 755 OR4XD1BWP7T $T=131440 474720 1 0 $X=131150 $Y=470510
X1908 107 104 103 768 2 1 770 OR4XD1BWP7T $T=149360 427680 1 180 $X=144590 $Y=427445
X1909 126 2 108 102 796 94 1 INR4D2BWP7T $T=156080 474720 0 180 $X=141230 $Y=470510
X1910 735 679 738 760 771 1 2 AO211D2BWP7T $T=140400 459040 1 0 $X=140110 $Y=454830
X1911 591 1 78 80 2 81 715 OAI211D0BWP7T $T=107920 419840 1 0 $X=107630 $Y=415630
X1912 515 1 596 83 2 10 716 OAI211D0BWP7T $T=114640 427680 0 180 $X=110990 $Y=423470
X1913 736 1 664 83 2 85 743 OAI211D0BWP7T $T=129760 427680 1 180 $X=126110 $Y=427445
X1914 718 1 724 733 2 744 748 OAI211D0BWP7T $T=128080 466880 0 0 $X=127790 $Y=466645
X1915 754 1 761 646 2 744 764 OAI211D0BWP7T $T=138720 466880 0 0 $X=138430 $Y=466645
X1916 475 1 589 592 2 CKND2D1BWP7T $T=69280 451200 1 0 $X=68990 $Y=446990
X1917 759 1 757 687 2 CKND2D1BWP7T $T=138160 451200 0 180 $X=135630 $Y=446990
X1918 742 1 758 87 2 CKND2D1BWP7T $T=140400 435520 0 180 $X=137870 $Y=431310
X1919 754 1 761 744 767 646 2 OAI211D2BWP7T $T=137600 466880 1 0 $X=137310 $Y=462670
X1920 523 1 659 678 2 CKND2D0BWP7T $T=100640 451200 0 0 $X=100350 $Y=450965
X1921 742 1 80 731 2 CKND2D0BWP7T $T=137600 419840 1 180 $X=135070 $Y=419605
X1922 84 1 708 728 2 CKND2D3BWP7T $T=140400 419840 0 180 $X=135070 $Y=415630
X1923 618 464 11 474 1 2 610 AO211D0BWP7T $T=84960 427680 1 180 $X=80750 $Y=427445
X1924 80 7 18 716 1 2 693 AO211D0BWP7T $T=115200 419840 1 180 $X=110990 $Y=419605
X1925 701 706 751 745 1 2 756 AO211D0BWP7T $T=133120 443360 0 0 $X=132830 $Y=443125
X1926 496 2 23 514 19 512 1 AOI211D2BWP7T $T=41280 427680 0 0 $X=40990 $Y=427445
X1927 619 2 623 654 464 66 1 AOI211D2BWP7T $T=91120 427680 1 0 $X=90830 $Y=423470
X1928 563 2 482 695 7 758 1 AOI211D2BWP7T $T=132000 443360 1 0 $X=131710 $Y=439150
X1929 4 2 11 458 1 NR2D3BWP7T $T=21120 443360 0 0 $X=20830 $Y=443125
X1930 3 2 471 8 1 NR2D3BWP7T $T=22240 474720 1 0 $X=21950 $Y=470510
X1931 15 2 482 12 1 NR2D3BWP7T $T=24480 419840 1 0 $X=24190 $Y=415630
X1932 458 2 483 16 1 NR2D3BWP7T $T=24480 451200 1 0 $X=24190 $Y=446990
X1933 17 2 481 13 1 NR2D3BWP7T $T=26160 459040 1 0 $X=25870 $Y=454830
X1934 466 2 536 483 1 NR2D3BWP7T $T=56400 435520 0 180 $X=51070 $Y=431310
X1935 722 2 495 742 1 NR2D3BWP7T $T=137040 435520 0 180 $X=131710 $Y=431310
X1936 660 735 1 2 705 751 744 MOAI22D0BWP7T $T=130320 451200 1 0 $X=130030 $Y=446990
X1937 48 521 1 2 50 AN2D1BWP7T $T=65360 427680 1 0 $X=65070 $Y=423470
X1938 37 575 1 2 585 AN2D1BWP7T $T=65920 419840 0 0 $X=65630 $Y=419605
X1939 84 512 1 2 32 AN2D1BWP7T $T=115200 419840 0 180 $X=112110 $Y=415630
X1940 747 742 1 2 480 AN2D1BWP7T $T=132000 419840 1 180 $X=128910 $Y=419605
X1941 512 10 86 1 2 ND2D2BWP7T $T=123040 419840 1 0 $X=122750 $Y=415630
X1942 710 2 676 706 706 1 671 724 AOI221D1BWP7T $T=110160 474720 1 0 $X=109870 $Y=470510
X1943 528 1 2 606 18 609 NR3D0BWP7T $T=79920 443360 1 0 $X=79630 $Y=439150
X1944 715 1 2 14 690 707 NR3D0BWP7T $T=110160 435520 1 0 $X=109870 $Y=431310
X1945 706 688 1 683 702 2 AOI21D1BWP7T $T=110160 474720 0 180 $X=106510 $Y=470510
X1946 51 50 490 549 2 1 ND3D2BWP7T $T=68160 427680 1 0 $X=67870 $Y=423470
X1947 56 673 553 492 2 1 ND3D2BWP7T $T=105120 474720 0 180 $X=99790 $Y=470510
X1948 641 2 67 659 1 NR2D0BWP7T $T=100080 435520 0 180 $X=97550 $Y=431310
X1949 465 468 477 22 485 1 2 ND4D2BWP7T $T=23920 459040 0 0 $X=23630 $Y=458805
X1950 486 531 30 544 534 1 2 ND4D2BWP7T $T=48560 474720 1 0 $X=48270 $Y=470510
X1951 498 57 633 497 595 1 2 ND4D2BWP7T $T=83840 427680 1 0 $X=83550 $Y=423470
X1952 608 1 617 605 490 595 2 OAI31D2BWP7T $T=81600 451200 1 0 $X=81310 $Y=446990
X1953 508 1 507 506 2 469 ND3D1BWP7T $T=46320 443360 0 180 $X=42670 $Y=439150
X1954 529 1 36 498 2 539 ND3D1BWP7T $T=51360 427680 0 0 $X=51070 $Y=427445
X1955 582 1 537 585 2 590 ND3D1BWP7T $T=66480 451200 0 0 $X=66190 $Y=450965
X1956 475 1 572 593 2 513 ND3D1BWP7T $T=68720 435520 1 0 $X=68430 $Y=431310
X1957 562 1 570 51 2 520 ND3D1BWP7T $T=68720 466880 1 0 $X=68430 $Y=462670
X1958 532 1 536 585 2 603 ND3D1BWP7T $T=69840 451200 0 0 $X=69550 $Y=450965
X1959 519 2 463 512 1 506 31 AOI211D1BWP7T $T=51360 427680 1 180 $X=47710 $Y=427445
X1960 528 1 473 507 516 494 2 IND4D2BWP7T $T=51920 443360 1 180 $X=43230 $Y=443125
X1961 22 2 502 472 1 INR2D1BWP7T $T=45760 427680 0 180 $X=42670 $Y=423470
.ENDS
***************************************
.SUBCKT ICV_17 1 2
** N=2 EP=2 IP=4 FDC=6
X1 1 2 DCAP8BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_18
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT CKBD2BWP7T I Z VDD VSS
** N=5 EP=4 IP=0 FDC=6
M0 VSS I 5 VSS N L=1.8e-07 W=5.25e-07 $X=1120 $Y=460 $D=0
M1 Z 5 VSS VSS N L=1.8e-07 W=5.25e-07 $X=1840 $Y=460 $D=0
M2 VSS 5 Z VSS N L=1.8e-07 W=5.25e-07 $X=2560 $Y=460 $D=0
M3 VDD I 5 VDD P L=1.8e-07 W=1.54e-06 $X=1120 $Y=2035 $D=16
M4 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1840 $Y=2205 $D=16
M5 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=2560 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AO221D0BWP7T B2 A1 A2 B1 C VSS VDD Z
** N=13 EP=8 IP=0 FDC=12
M0 11 A1 9 VSS N L=1.8e-07 W=5e-07 $X=1075 $Y=775 $D=0
M1 VSS A2 11 VSS N L=1.8e-07 W=5e-07 $X=1520 $Y=775 $D=0
M2 12 B2 VSS VSS N L=1.8e-07 W=5e-07 $X=2290 $Y=520 $D=0
M3 9 B1 12 VSS N L=1.8e-07 W=5e-07 $X=2720 $Y=520 $D=0
M4 VSS C 9 VSS N L=1.8e-07 W=5e-07 $X=3440 $Y=520 $D=0
M5 Z 9 VSS VSS N L=1.8e-07 W=5e-07 $X=4240 $Y=520 $D=0
M6 13 B2 10 VDD P L=1.8e-07 W=6.85e-07 $X=640 $Y=2555 $D=16
M7 9 A1 13 VDD P L=1.8e-07 W=6.85e-07 $X=1360 $Y=2555 $D=16
M8 13 A2 9 VDD P L=1.8e-07 W=6.85e-07 $X=2080 $Y=2555 $D=16
M9 10 B1 13 VDD P L=1.8e-07 W=6.85e-07 $X=2800 $Y=2555 $D=16
M10 VDD C 10 VDD P L=1.8e-07 W=6.85e-07 $X=3520 $Y=2555 $D=16
M11 Z 9 VDD VDD P L=1.8e-07 W=6.85e-07 $X=4240 $Y=2555 $D=16
.ENDS
***************************************
.SUBCKT ICV_19 1 2
** N=2 EP=2 IP=4 FDC=8
X0 1 2 DCAP8BWP7T $T=0 0 0 0 $X=-290 $Y=-235
X1 2 1 DCAPBWP7T $T=4480 0 0 0 $X=4190 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_20
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21 1 2
** N=2 EP=2 IP=4 FDC=10
X0 1 2 ICV_3 $T=4480 0 0 0 $X=4190 $Y=-235
X1 1 2 DCAP8BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT FILL32BWP7T
** N=35 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DFCND1BWP7T CP D CDN QN VDD VSS Q
** N=20 EP=7 IP=0 FDC=30
M0 VSS CP 8 VSS N L=1.8e-07 W=5e-07 $X=640 $Y=840 $D=0
M1 9 8 VSS VSS N L=1.8e-07 W=5e-07 $X=1240 $Y=840 $D=0
M2 16 8 VSS VSS N L=1.8e-07 W=9.4e-07 $X=2660 $Y=405 $D=0
M3 11 D 16 VSS N L=1.8e-07 W=9.4e-07 $X=3160 $Y=405 $D=0
M4 17 9 11 VSS N L=1.8e-07 W=4.2e-07 $X=4005 $Y=895 $D=0
M5 18 CDN 17 VSS N L=1.8e-07 W=4.2e-07 $X=4435 $Y=895 $D=0
M6 VSS 12 18 VSS N L=1.8e-07 W=4.2e-07 $X=4865 $Y=895 $D=0
M7 12 11 VSS VSS N L=1.8e-07 W=5.4e-07 $X=5715 $Y=775 $D=0
M8 14 9 12 VSS N L=1.8e-07 W=9.1e-07 $X=6435 $Y=405 $D=0
M9 13 8 14 VSS N L=1.8e-07 W=4.2e-07 $X=7155 $Y=895 $D=0
M10 VSS 15 13 VSS N L=1.8e-07 W=4.2e-07 $X=8730 $Y=895 $D=0
M11 19 CDN VSS VSS N L=1.8e-07 W=9.7e-07 $X=9330 $Y=345 $D=0
M12 15 14 19 VSS N L=1.8e-07 W=9.7e-07 $X=9760 $Y=345 $D=0
M13 VSS 13 QN VSS N L=1.8e-07 W=9.4e-07 $X=11360 $Y=405 $D=0
M14 Q 15 VSS VSS N L=1.8e-07 W=1e-06 $X=12080 $Y=345 $D=0
M15 VDD CP 8 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2345 $D=16
M16 9 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1240 $Y=2345 $D=16
M17 20 9 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2525 $Y=2205 $D=16
M18 11 D 20 VDD P L=1.8e-07 W=1.37e-06 $X=2955 $Y=2205 $D=16
M19 10 8 11 VDD P L=1.8e-07 W=4.2e-07 $X=3795 $Y=2365 $D=16
M20 VDD CDN 10 VDD P L=1.8e-07 W=4.2e-07 $X=4515 $Y=2365 $D=16
M21 10 12 VDD VDD P L=1.8e-07 W=4.2e-07 $X=5115 $Y=2365 $D=16
M22 12 11 VDD VDD P L=1.8e-07 W=6.2e-07 $X=6375 $Y=2175 $D=16
M23 14 8 12 VDD P L=1.8e-07 W=6.2e-07 $X=7255 $Y=2175 $D=16
M24 13 9 14 VDD P L=1.8e-07 W=4.2e-07 $X=8070 $Y=2175 $D=16
M25 VDD 15 13 VDD P L=1.8e-07 W=6e-07 $X=8790 $Y=2175 $D=16
M26 15 CDN VDD VDD P L=1.8e-07 W=4.2e-07 $X=9390 $Y=3095 $D=16
M27 VDD 14 15 VDD P L=1.8e-07 W=1.37e-06 $X=10150 $Y=2205 $D=16
M28 VDD 13 QN VDD P L=1.8e-07 W=8.35e-07 $X=11410 $Y=2205 $D=16
M29 Q 15 VDD VDD P L=1.8e-07 W=1.37e-06 $X=12080 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT XNR2D2BWP7T A1 A2 ZN VSS VDD
** N=9 EP=5 IP=0 FDC=14
M0 VSS 8 7 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 6 A1 VSS VSS N L=1.8e-07 W=5e-07 $X=1380 $Y=845 $D=0
M2 9 6 7 VSS N L=1.8e-07 W=5e-07 $X=2960 $Y=845 $D=0
M3 8 A1 9 VSS N L=1.8e-07 W=5e-07 $X=3680 $Y=845 $D=0
M4 VSS A2 8 VSS N L=1.8e-07 W=1e-06 $X=4400 $Y=345 $D=0
M5 ZN 9 VSS VSS N L=1.8e-07 W=1e-06 $X=5200 $Y=345 $D=0
M6 VSS 9 ZN VSS N L=1.8e-07 W=1e-06 $X=5920 $Y=345 $D=0
M7 VDD 8 7 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M8 6 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1420 $Y=2205 $D=16
M9 9 A1 7 VDD P L=1.8e-07 W=6.85e-07 $X=2960 $Y=2595 $D=16
M10 8 6 9 VDD P L=1.8e-07 W=6.85e-07 $X=3735 $Y=2205 $D=16
M11 VDD A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=4455 $Y=2205 $D=16
M12 ZN 9 VDD VDD P L=1.8e-07 W=1.37e-06 $X=5200 $Y=2205 $D=16
M13 VDD 9 ZN VDD P L=1.8e-07 W=1.37e-06 $X=5920 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AOI211XD0BWP7T C VSS VDD B A2 ZN A1
** N=10 EP=7 IP=0 FDC=8
M0 ZN C VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=680 $D=0
M1 VSS B ZN VSS N L=1.8e-07 W=5e-07 $X=1340 $Y=680 $D=0
M2 9 A2 VSS VSS N L=1.8e-07 W=5e-07 $X=2060 $Y=680 $D=0
M3 ZN A1 9 VSS N L=1.8e-07 W=5e-07 $X=2560 $Y=680 $D=0
M4 10 C VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M5 8 B 10 VDD P L=1.8e-07 W=1.37e-06 $X=1100 $Y=2205 $D=16
M6 ZN A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=1830 $Y=2205 $D=16
M7 8 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2560 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT DFCND2BWP7T CP D CDN QN Q VSS VDD
** N=20 EP=7 IP=0 FDC=34
M0 VSS CP 8 VSS N L=1.8e-07 W=5e-07 $X=640 $Y=840 $D=0
M1 9 8 VSS VSS N L=1.8e-07 W=5e-07 $X=1240 $Y=840 $D=0
M2 16 8 VSS VSS N L=1.8e-07 W=9.4e-07 $X=2660 $Y=405 $D=0
M3 11 D 16 VSS N L=1.8e-07 W=9.4e-07 $X=3160 $Y=405 $D=0
M4 17 9 11 VSS N L=1.8e-07 W=4.2e-07 $X=4005 $Y=895 $D=0
M5 18 CDN 17 VSS N L=1.8e-07 W=4.2e-07 $X=4435 $Y=895 $D=0
M6 VSS 12 18 VSS N L=1.8e-07 W=4.2e-07 $X=4865 $Y=895 $D=0
M7 12 11 VSS VSS N L=1.8e-07 W=5.4e-07 $X=5715 $Y=775 $D=0
M8 13 9 12 VSS N L=1.8e-07 W=9.1e-07 $X=6435 $Y=405 $D=0
M9 14 8 13 VSS N L=1.8e-07 W=4.2e-07 $X=7155 $Y=895 $D=0
M10 VSS 15 14 VSS N L=1.8e-07 W=9.7e-07 $X=8870 $Y=345 $D=0
M11 19 CDN VSS VSS N L=1.8e-07 W=9.7e-07 $X=9670 $Y=345 $D=0
M12 15 13 19 VSS N L=1.8e-07 W=9.7e-07 $X=10100 $Y=345 $D=0
M13 QN 14 VSS VSS N L=1.8e-07 W=1e-06 $X=11600 $Y=345 $D=0
M14 VSS 14 QN VSS N L=1.8e-07 W=1e-06 $X=12320 $Y=345 $D=0
M15 Q 15 VSS VSS N L=1.8e-07 W=1e-06 $X=13040 $Y=345 $D=0
M16 VSS 15 Q VSS N L=1.8e-07 W=1e-06 $X=13760 $Y=345 $D=0
M17 VDD CP 8 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2345 $D=16
M18 9 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1240 $Y=2345 $D=16
M19 20 9 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2525 $Y=2205 $D=16
M20 11 D 20 VDD P L=1.8e-07 W=1.37e-06 $X=2955 $Y=2205 $D=16
M21 10 8 11 VDD P L=1.8e-07 W=4.2e-07 $X=3795 $Y=2365 $D=16
M22 VDD CDN 10 VDD P L=1.8e-07 W=4.2e-07 $X=4515 $Y=2365 $D=16
M23 10 12 VDD VDD P L=1.8e-07 W=4.2e-07 $X=5115 $Y=2365 $D=16
M24 12 11 VDD VDD P L=1.8e-07 W=6.2e-07 $X=6375 $Y=2175 $D=16
M25 13 8 12 VDD P L=1.8e-07 W=6.2e-07 $X=7255 $Y=2175 $D=16
M26 14 9 13 VDD P L=1.8e-07 W=4.2e-07 $X=8070 $Y=2175 $D=16
M27 VDD 15 14 VDD P L=1.8e-07 W=9.7e-07 $X=9010 $Y=2175 $D=16
M28 15 CDN VDD VDD P L=1.8e-07 W=4.2e-07 $X=9850 $Y=3095 $D=16
M29 VDD 13 15 VDD P L=1.8e-07 W=1.23e-06 $X=10620 $Y=2345 $D=16
M30 QN 14 VDD VDD P L=1.8e-07 W=1.23e-06 $X=11560 $Y=2345 $D=16
M31 VDD 14 QN VDD P L=1.8e-07 W=1.37e-06 $X=12320 $Y=2205 $D=16
M32 Q 15 VDD VDD P L=1.8e-07 W=1.37e-06 $X=13040 $Y=2205 $D=16
M33 VDD 15 Q VDD P L=1.8e-07 W=1.37e-06 $X=13760 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OAI21D2BWP7T B VSS ZN A1 A2 VDD
** N=9 EP=6 IP=0 FDC=12
M0 VSS B 7 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 7 B VSS VSS N L=1.8e-07 W=1e-06 $X=1345 $Y=345 $D=0
M2 ZN A2 7 VSS N L=1.8e-07 W=1e-06 $X=2080 $Y=345 $D=0
M3 7 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=2800 $Y=345 $D=0
M4 ZN A1 7 VSS N L=1.8e-07 W=1e-06 $X=3520 $Y=345 $D=0
M5 7 A2 ZN VSS N L=1.8e-07 W=1e-06 $X=4240 $Y=345 $D=0
M6 ZN B VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M7 VDD B ZN VDD P L=1.8e-07 W=1.37e-06 $X=1345 $Y=2205 $D=16
M8 8 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2145 $Y=2205 $D=16
M9 ZN A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=2800 $Y=2205 $D=16
M10 9 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3520 $Y=2205 $D=16
M11 VDD A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=4200 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IOA21D1BWP7T A1 A2 VSS ZN B VDD
** N=9 EP=6 IP=0 FDC=8
M0 8 A1 7 VSS N L=1.8e-07 W=5e-07 $X=625 $Y=345 $D=0
M1 VSS A2 8 VSS N L=1.8e-07 W=5e-07 $X=1205 $Y=345 $D=0
M2 9 7 VSS VSS N L=1.8e-07 W=1e-06 $X=1975 $Y=345 $D=0
M3 ZN B 9 VSS N L=1.8e-07 W=1e-06 $X=2560 $Y=345 $D=0
M4 7 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=465 $Y=2205 $D=16
M5 VDD A2 7 VDD P L=1.8e-07 W=6.85e-07 $X=1185 $Y=2205 $D=16
M6 ZN 7 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1840 $Y=2205 $D=16
M7 VDD B ZN VDD P L=1.8e-07 W=1.37e-06 $X=2560 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OAI22D1BWP7T B1 B2 VSS A2 VDD ZN A1
** N=10 EP=7 IP=0 FDC=8
M0 VSS B1 8 VSS N L=1.8e-07 W=1e-06 $X=640 $Y=345 $D=0
M1 8 B2 VSS VSS N L=1.8e-07 W=1e-06 $X=1440 $Y=345 $D=0
M2 ZN A2 8 VSS N L=1.8e-07 W=1e-06 $X=2180 $Y=345 $D=0
M3 8 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=3120 $Y=345 $D=0
M4 9 B1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=640 $Y=2205 $D=16
M5 VDD B2 9 VDD P L=1.8e-07 W=1.37e-06 $X=1440 $Y=2205 $D=16
M6 10 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2420 $Y=2205 $D=16
M7 ZN A1 10 VDD P L=1.8e-07 W=1.37e-06 $X=3120 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT DEL1BWP7T I VSS VDD Z
** N=7 EP=4 IP=0 FDC=8
M0 VSS I 5 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=515 $D=0
M1 6 5 VSS VSS N L=7e-07 W=8.3e-07 $X=1340 $Y=515 $D=0
M2 VSS 6 7 VSS N L=7e-07 W=6e-07 $X=3520 $Y=505 $D=0
M3 Z 7 VSS VSS N L=1.8e-07 W=1e-06 $X=4760 $Y=345 $D=0
M4 VDD I 5 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2795 $D=16
M5 6 5 VDD VDD P L=7e-07 W=1.2e-06 $X=1340 $Y=2280 $D=16
M6 VDD 6 7 VDD P L=7e-07 W=9e-07 $X=3520 $Y=2675 $D=16
M7 Z 7 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4760 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AO221D1BWP7T A2 A1 B2 B1 C VSS VDD Z
** N=13 EP=8 IP=0 FDC=12
M0 12 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 11 A1 12 VSS N L=1.8e-07 W=1e-06 $X=1260 $Y=345 $D=0
M2 13 B2 VSS VSS N L=1.8e-07 W=1e-06 $X=2685 $Y=345 $D=0
M3 11 B1 13 VSS N L=1.8e-07 W=1e-06 $X=3230 $Y=345 $D=0
M4 VSS C 11 VSS N L=1.8e-07 W=1e-06 $X=4065 $Y=345 $D=0
M5 Z 11 VSS VSS N L=1.8e-07 W=1e-06 $X=4800 $Y=345 $D=0
M6 11 A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M7 9 A1 11 VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M8 9 B2 10 VDD P L=1.8e-07 W=1.37e-06 $X=2640 $Y=2205 $D=16
M9 10 B1 9 VDD P L=1.8e-07 W=1.37e-06 $X=3360 $Y=2205 $D=16
M10 VDD C 10 VDD P L=1.8e-07 W=1.37e-06 $X=4080 $Y=2205 $D=16
M11 Z 11 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4800 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT DFCND0BWP7T CP D CDN QN VDD VSS Q
** N=20 EP=7 IP=0 FDC=30
M0 VSS CP 8 VSS N L=1.8e-07 W=5e-07 $X=640 $Y=840 $D=0
M1 9 8 VSS VSS N L=1.8e-07 W=5e-07 $X=1240 $Y=840 $D=0
M2 16 8 VSS VSS N L=1.8e-07 W=9.4e-07 $X=2660 $Y=405 $D=0
M3 11 D 16 VSS N L=1.8e-07 W=9.4e-07 $X=3160 $Y=405 $D=0
M4 17 9 11 VSS N L=1.8e-07 W=4.2e-07 $X=4005 $Y=895 $D=0
M5 18 CDN 17 VSS N L=1.8e-07 W=4.2e-07 $X=4435 $Y=895 $D=0
M6 VSS 12 18 VSS N L=1.8e-07 W=4.2e-07 $X=4865 $Y=895 $D=0
M7 12 11 VSS VSS N L=1.8e-07 W=5.4e-07 $X=5715 $Y=775 $D=0
M8 14 9 12 VSS N L=1.8e-07 W=9.1e-07 $X=6435 $Y=405 $D=0
M9 13 8 14 VSS N L=1.8e-07 W=4.2e-07 $X=7155 $Y=895 $D=0
M10 VSS 15 13 VSS N L=1.8e-07 W=4.2e-07 $X=8730 $Y=895 $D=0
M11 19 CDN VSS VSS N L=1.8e-07 W=9.7e-07 $X=9330 $Y=345 $D=0
M12 15 14 19 VSS N L=1.8e-07 W=9.7e-07 $X=9760 $Y=345 $D=0
M13 VSS 13 QN VSS N L=1.8e-07 W=5e-07 $X=11360 $Y=540 $D=0
M14 Q 15 VSS VSS N L=1.8e-07 W=5e-07 $X=12080 $Y=540 $D=0
M15 VDD CP 8 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2345 $D=16
M16 9 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1240 $Y=2345 $D=16
M17 20 9 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2525 $Y=2205 $D=16
M18 11 D 20 VDD P L=1.8e-07 W=1.37e-06 $X=2955 $Y=2205 $D=16
M19 10 8 11 VDD P L=1.8e-07 W=4.2e-07 $X=3795 $Y=2365 $D=16
M20 VDD CDN 10 VDD P L=1.8e-07 W=4.2e-07 $X=4515 $Y=2365 $D=16
M21 10 12 VDD VDD P L=1.8e-07 W=4.2e-07 $X=5115 $Y=2365 $D=16
M22 12 11 VDD VDD P L=1.8e-07 W=6.2e-07 $X=6375 $Y=2175 $D=16
M23 14 8 12 VDD P L=1.8e-07 W=6.2e-07 $X=7255 $Y=2175 $D=16
M24 13 9 14 VDD P L=1.8e-07 W=4.2e-07 $X=8070 $Y=2175 $D=16
M25 VDD 15 13 VDD P L=1.8e-07 W=6e-07 $X=8790 $Y=2175 $D=16
M26 15 CDN VDD VDD P L=1.8e-07 W=4.2e-07 $X=9390 $Y=3095 $D=16
M27 VDD 14 15 VDD P L=1.8e-07 W=1.31e-06 $X=10150 $Y=2205 $D=16
M28 VDD 13 QN VDD P L=1.8e-07 W=6.85e-07 $X=11410 $Y=2205 $D=16
M29 Q 15 VDD VDD P L=1.8e-07 W=6.85e-07 $X=12080 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OA222D0BWP7T C1 C2 B2 A2 A1 B1 VDD Z VSS
** N=15 EP=9 IP=0 FDC=14
M0 VSS C1 10 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=565 $D=0
M1 10 C2 VSS VSS N L=1.8e-07 W=5e-07 $X=1340 $Y=565 $D=0
M2 12 B2 10 VSS N L=1.8e-07 W=5e-07 $X=2060 $Y=565 $D=0
M3 11 A2 12 VSS N L=1.8e-07 W=5e-07 $X=2660 $Y=780 $D=0
M4 12 A1 11 VSS N L=1.8e-07 W=5e-07 $X=3380 $Y=780 $D=0
M5 10 B1 12 VSS N L=1.8e-07 W=5e-07 $X=3980 $Y=360 $D=0
M6 Z 11 VSS VSS N L=1.8e-07 W=5e-07 $X=5360 $Y=845 $D=0
M7 13 C1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2890 $D=16
M8 11 C2 13 VDD P L=1.8e-07 W=6.85e-07 $X=1220 $Y=2890 $D=16
M9 14 B2 11 VDD P L=1.8e-07 W=6.85e-07 $X=1995 $Y=2890 $D=16
M10 VDD B1 14 VDD P L=1.8e-07 W=6.85e-07 $X=2490 $Y=2890 $D=16
M11 15 A2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=3295 $Y=2890 $D=16
M12 11 A1 15 VDD P L=1.8e-07 W=6.85e-07 $X=3900 $Y=2890 $D=16
M13 Z 11 VDD VDD P L=1.8e-07 W=6.85e-07 $X=5360 $Y=2890 $D=16
.ENDS
***************************************
.SUBCKT AOI211XD1BWP7T C VDD B VSS ZN A1 A2
** N=10 EP=7 IP=0 FDC=12
M0 ZN C VSS VSS N L=1.8e-07 W=1e-06 $X=1730 $Y=345 $D=0
M1 VSS B ZN VSS N L=1.8e-07 W=1e-06 $X=2860 $Y=345 $D=0
M2 10 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=3820 $Y=345 $D=0
M3 ZN A1 10 VSS N L=1.8e-07 W=1e-06 $X=4555 $Y=345 $D=0
M4 8 B 9 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M5 VDD C 8 VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M6 8 C VDD VDD P L=1.8e-07 W=1.37e-06 $X=2140 $Y=2205 $D=16
M7 9 B 8 VDD P L=1.8e-07 W=1.37e-06 $X=2860 $Y=2205 $D=16
M8 ZN A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=3580 $Y=2205 $D=16
M9 9 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4360 $Y=2205 $D=16
M10 ZN A1 9 VDD P L=1.8e-07 W=1.37e-06 $X=5160 $Y=2205 $D=16
M11 9 A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=5885 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INVD2P5BWP7T I ZN VSS VDD
** N=4 EP=4 IP=0 FDC=6
M0 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 VSS I ZN VSS N L=1.8e-07 W=4.65e-07 $X=2060 $Y=880 $D=0
M3 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M4 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M5 VDD I ZN VDD P L=1.8e-07 W=6.85e-07 $X=2060 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INVD6BWP7T I ZN VSS VDD
** N=4 EP=4 IP=0 FDC=12
M0 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=2060 $Y=345 $D=0
M3 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=2780 $Y=345 $D=0
M4 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=3500 $Y=345 $D=0
M5 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=4220 $Y=345 $D=0
M6 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M7 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M8 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M9 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M10 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=3500 $Y=2205 $D=16
M11 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=4220 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OAI222D2BWP7T C2 C1 VSS B2 B1 A1 A2 VDD ZN
** N=17 EP=9 IP=0 FDC=24
M0 VSS C1 10 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 10 C2 VSS VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 VSS C2 10 VSS N L=1.8e-07 W=1e-06 $X=2060 $Y=345 $D=0
M3 10 C1 VSS VSS N L=1.8e-07 W=1e-06 $X=2780 $Y=345 $D=0
M4 11 B1 10 VSS N L=1.8e-07 W=1e-06 $X=3500 $Y=345 $D=0
M5 10 B2 11 VSS N L=1.8e-07 W=1e-06 $X=4220 $Y=345 $D=0
M6 11 B2 10 VSS N L=1.8e-07 W=1e-06 $X=4940 $Y=345 $D=0
M7 10 B1 11 VSS N L=1.8e-07 W=1e-06 $X=5660 $Y=345 $D=0
M8 11 A2 ZN VSS N L=1.8e-07 W=1e-06 $X=7080 $Y=345 $D=0
M9 ZN A1 11 VSS N L=1.8e-07 W=1e-06 $X=7800 $Y=345 $D=0
M10 11 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=8520 $Y=345 $D=0
M11 ZN A2 11 VSS N L=1.8e-07 W=1e-06 $X=9240 $Y=345 $D=0
M12 12 C1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M13 ZN C2 12 VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M14 13 C2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M15 VDD C1 13 VDD P L=1.8e-07 W=1.37e-06 $X=2560 $Y=2205 $D=16
M16 14 B1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3440 $Y=2205 $D=16
M17 ZN B2 14 VDD P L=1.8e-07 W=1.37e-06 $X=4220 $Y=2205 $D=16
M18 15 B2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4940 $Y=2205 $D=16
M19 VDD B1 15 VDD P L=1.8e-07 W=1.37e-06 $X=5520 $Y=2205 $D=16
M20 16 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=7080 $Y=2205 $D=16
M21 ZN A1 16 VDD P L=1.8e-07 W=1.37e-06 $X=7800 $Y=2205 $D=16
M22 17 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=8520 $Y=2205 $D=16
M23 VDD A2 17 VDD P L=1.8e-07 W=1.37e-06 $X=9040 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INVD5BWP7T I VSS VDD ZN
** N=4 EP=4 IP=0 FDC=10
M0 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=720 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=1440 $Y=345 $D=0
M2 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=2200 $Y=345 $D=0
M3 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=2920 $Y=345 $D=0
M4 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=3680 $Y=345 $D=0
M5 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=720 $Y=2205 $D=16
M6 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1440 $Y=2205 $D=16
M7 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=2200 $Y=2205 $D=16
M8 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=2920 $Y=2205 $D=16
M9 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=3680 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT XOR2D2BWP7T A1 A2 Z VSS VDD
** N=9 EP=5 IP=0 FDC=14
M0 VSS 8 7 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 6 A1 VSS VSS N L=1.8e-07 W=5e-07 $X=1425 $Y=845 $D=0
M2 9 A1 7 VSS N L=1.8e-07 W=8.1e-07 $X=2970 $Y=535 $D=0
M3 8 6 9 VSS N L=1.8e-07 W=8.1e-07 $X=3730 $Y=535 $D=0
M4 VSS A2 8 VSS N L=1.8e-07 W=1e-06 $X=4450 $Y=345 $D=0
M5 Z 9 VSS VSS N L=1.8e-07 W=1e-06 $X=5170 $Y=345 $D=0
M6 VSS 9 Z VSS N L=1.8e-07 W=1e-06 $X=5890 $Y=345 $D=0
M7 VDD 8 7 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M8 6 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1425 $Y=2205 $D=16
M9 9 6 7 VDD P L=1.8e-07 W=7.3e-07 $X=2960 $Y=2320 $D=16
M10 8 A1 9 VDD P L=1.8e-07 W=7.3e-07 $X=3680 $Y=2635 $D=16
M11 VDD A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=4450 $Y=2205 $D=16
M12 Z 9 VDD VDD P L=1.8e-07 W=1.37e-06 $X=5170 $Y=2205 $D=16
M13 VDD 9 Z VDD P L=1.8e-07 W=1.37e-06 $X=5890 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR2D2P5BWP7T A2 VDD VSS A1 ZN
** N=8 EP=5 IP=0 FDC=12
M0 ZN A2 VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS A1 ZN VSS N L=1.8e-07 W=1e-06 $X=1350 $Y=345 $D=0
M2 ZN A1 VSS VSS N L=1.8e-07 W=1e-06 $X=2110 $Y=345 $D=0
M3 VSS A2 ZN VSS N L=1.8e-07 W=1e-06 $X=2830 $Y=345 $D=0
M4 ZN A2 VSS VSS N L=1.8e-07 W=5e-07 $X=3590 $Y=845 $D=0
M5 VSS A1 ZN VSS N L=1.8e-07 W=5e-07 $X=4350 $Y=845 $D=0
M6 6 A2 VDD VDD P L=1.8e-07 W=1.14e-06 $X=620 $Y=2435 $D=16
M7 ZN A1 6 VDD P L=1.8e-07 W=1.14e-06 $X=1220 $Y=2435 $D=16
M8 7 A1 ZN VDD P L=1.8e-07 W=1.14e-06 $X=1940 $Y=2435 $D=16
M9 VDD A2 7 VDD P L=1.8e-07 W=1.14e-06 $X=2660 $Y=2435 $D=16
M10 8 A2 VDD VDD P L=1.8e-07 W=1.14e-06 $X=3380 $Y=2435 $D=16
M11 ZN A1 8 VDD P L=1.8e-07 W=1.14e-06 $X=4150 $Y=2435 $D=16
.ENDS
***************************************
.SUBCKT OAI31D0BWP7T A1 A2 A3 ZN B VSS VDD
** N=10 EP=7 IP=0 FDC=8
M0 8 A1 ZN VSS N L=1.8e-07 W=5e-07 $X=620 $Y=845 $D=0
M1 ZN A2 8 VSS N L=1.8e-07 W=5e-07 $X=1220 $Y=845 $D=0
M2 8 A3 ZN VSS N L=1.8e-07 W=5e-07 $X=1945 $Y=845 $D=0
M3 VSS B 8 VSS N L=1.8e-07 W=5e-07 $X=2560 $Y=845 $D=0
M4 9 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2755 $D=16
M5 10 A2 9 VDD P L=1.8e-07 W=6.85e-07 $X=1210 $Y=2755 $D=16
M6 ZN A3 10 VDD P L=1.8e-07 W=6.85e-07 $X=1800 $Y=2755 $D=16
M7 VDD B ZN VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2755 $D=16
.ENDS
***************************************
.SUBCKT CKAN2D2BWP7T A1 A2 Z VDD VSS
** N=7 EP=5 IP=0 FDC=8
M0 7 A1 6 VSS N L=1.8e-07 W=7.4e-07 $X=705 $Y=345 $D=0
M1 VSS A2 7 VSS N L=1.8e-07 W=7.4e-07 $X=1480 $Y=345 $D=0
M2 Z 6 VSS VSS N L=1.8e-07 W=5.25e-07 $X=2400 $Y=345 $D=0
M3 VSS 6 Z VSS N L=1.8e-07 W=5.25e-07 $X=3120 $Y=345 $D=0
M4 6 A1 VDD VDD P L=1.8e-07 W=1.23e-06 $X=705 $Y=2345 $D=16
M5 VDD A2 6 VDD P L=1.8e-07 W=1.29e-06 $X=1480 $Y=2285 $D=16
M6 Z 6 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2400 $Y=2205 $D=16
M7 VDD 6 Z VDD P L=1.8e-07 W=1.37e-06 $X=3120 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKAN2D1BWP7T A1 A2 VSS VDD Z
** N=7 EP=5 IP=0 FDC=6
M0 7 A1 6 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=515 $D=0
M1 VSS A2 7 VSS N L=1.8e-07 W=5e-07 $X=1090 $Y=515 $D=0
M2 Z 6 VSS VSS N L=1.8e-07 W=5.25e-07 $X=2000 $Y=515 $D=0
M3 6 A1 VDD VDD P L=1.8e-07 W=8.5e-07 $X=520 $Y=2205 $D=16
M4 VDD A2 6 VDD P L=1.8e-07 W=9e-07 $X=1240 $Y=2205 $D=16
M5 Z 6 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2000 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKND4BWP7T I ZN VSS VDD
** N=4 EP=4 IP=0 FDC=8
M0 VSS I ZN VSS N L=1.8e-07 W=7e-07 $X=1420 $Y=345 $D=0
M1 ZN I VSS VSS N L=1.8e-07 W=7e-07 $X=2140 $Y=345 $D=0
M2 VSS I ZN VSS N L=1.8e-07 W=7e-07 $X=2940 $Y=345 $D=0
M3 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=700 $Y=2205 $D=16
M4 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1420 $Y=2205 $D=16
M5 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=2220 $Y=2205 $D=16
M6 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=2940 $Y=2205 $D=16
D7 VSS I DN AREA=2.037e-13 PJ=1.81e-06 $X=140 $Y=860 $D=32
.ENDS
***************************************
.SUBCKT AN4D0BWP7T A1 A2 A3 A4 VDD VSS Z
** N=11 EP=7 IP=0 FDC=10
M0 9 A1 8 VSS N L=1.8e-07 W=5e-07 $X=625 $Y=345 $D=0
M1 10 A2 9 VSS N L=1.8e-07 W=5e-07 $X=1205 $Y=345 $D=0
M2 11 A3 10 VSS N L=1.8e-07 W=5e-07 $X=1785 $Y=345 $D=0
M3 VSS A4 11 VSS N L=1.8e-07 W=5e-07 $X=2365 $Y=345 $D=0
M4 Z 8 VSS VSS N L=1.8e-07 W=5e-07 $X=3105 $Y=345 $D=0
M5 8 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=460 $Y=2205 $D=16
M6 VDD A2 8 VDD P L=1.8e-07 W=6.85e-07 $X=1185 $Y=2205 $D=16
M7 8 A3 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1785 $Y=2205 $D=16
M8 VDD A4 8 VDD P L=1.8e-07 W=6.85e-07 $X=2515 $Y=2205 $D=16
M9 Z 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=3115 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR3D2BWP7T A3 VDD A2 A1 ZN VSS
** N=8 EP=6 IP=0 FDC=24
M0 ZN A3 VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=345 $D=0
M1 VSS A3 ZN VSS N L=1.8e-07 W=5e-07 $X=1340 $Y=345 $D=0
M2 ZN A3 VSS VSS N L=1.8e-07 W=5e-07 $X=2060 $Y=345 $D=0
M3 VSS A3 ZN VSS N L=1.8e-07 W=5e-07 $X=2780 $Y=345 $D=0
M4 ZN A2 VSS VSS N L=1.8e-07 W=5e-07 $X=3500 $Y=345 $D=0
M5 VSS A2 ZN VSS N L=1.8e-07 W=5e-07 $X=4220 $Y=345 $D=0
M6 ZN A2 VSS VSS N L=1.8e-07 W=5e-07 $X=4940 $Y=345 $D=0
M7 VSS A2 ZN VSS N L=1.8e-07 W=5e-07 $X=5660 $Y=345 $D=0
M8 ZN A1 VSS VSS N L=1.8e-07 W=5e-07 $X=7100 $Y=345 $D=0
M9 VSS A1 ZN VSS N L=1.8e-07 W=5e-07 $X=7820 $Y=345 $D=0
M10 ZN A1 VSS VSS N L=1.8e-07 W=5e-07 $X=8540 $Y=345 $D=0
M11 VSS A1 ZN VSS N L=1.8e-07 W=5e-07 $X=9260 $Y=345 $D=0
M12 VDD A3 7 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M13 7 A3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M14 VDD A3 7 VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M15 7 A3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M16 8 A2 7 VDD P L=1.8e-07 W=1.37e-06 $X=3500 $Y=2205 $D=16
M17 7 A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=4220 $Y=2205 $D=16
M18 8 A2 7 VDD P L=1.8e-07 W=1.37e-06 $X=4940 $Y=2205 $D=16
M19 7 A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=5660 $Y=2205 $D=16
M20 8 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=7100 $Y=2205 $D=16
M21 ZN A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=7820 $Y=2205 $D=16
M22 8 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=8540 $Y=2205 $D=16
M23 ZN A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=9260 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OR2D2BWP7T A1 A2 Z VSS VDD
** N=7 EP=5 IP=0 FDC=8
M0 6 A1 VSS VSS N L=1.8e-07 W=5e-07 $X=660 $Y=345 $D=0
M1 VSS A2 6 VSS N L=1.8e-07 W=5e-07 $X=1380 $Y=345 $D=0
M2 Z 6 VSS VSS N L=1.8e-07 W=1e-06 $X=2100 $Y=345 $D=0
M3 VSS 6 Z VSS N L=1.8e-07 W=1e-06 $X=2820 $Y=345 $D=0
M4 7 A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M5 VDD A2 7 VDD P L=1.8e-07 W=1.37e-06 $X=1380 $Y=2205 $D=16
M6 Z 6 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2200 $Y=2205 $D=16
M7 VDD 6 Z VDD P L=1.8e-07 W=1.37e-06 $X=2920 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IAO21D2BWP7T A1 A2 B ZN VDD VSS
** N=10 EP=6 IP=0 FDC=12
M0 7 A1 VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS A2 7 VSS N L=1.8e-07 W=1e-06 $X=1345 $Y=345 $D=0
M2 ZN 7 VSS VSS N L=1.8e-07 W=1e-06 $X=2065 $Y=345 $D=0
M3 VSS B ZN VSS N L=1.8e-07 W=1e-06 $X=2785 $Y=345 $D=0
M4 ZN B VSS VSS N L=1.8e-07 W=1e-06 $X=3505 $Y=345 $D=0
M5 VSS 7 ZN VSS N L=1.8e-07 W=1e-06 $X=4225 $Y=345 $D=0
M6 8 A1 7 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M7 VDD A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=1225 $Y=2205 $D=16
M8 9 7 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2125 $Y=2205 $D=16
M9 ZN B 9 VDD P L=1.8e-07 W=1.37e-06 $X=2785 $Y=2205 $D=16
M10 10 B ZN VDD P L=1.8e-07 W=1.37e-06 $X=3505 $Y=2205 $D=16
M11 VDD 7 10 VDD P L=1.8e-07 W=1.37e-06 $X=4225 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ND2D1P5BWP7T A1 ZN A2 VSS VDD
** N=7 EP=5 IP=0 FDC=8
M0 6 A2 VSS VSS N L=1.8e-07 W=7.5e-07 $X=740 $Y=345 $D=0
M1 ZN A1 6 VSS N L=1.8e-07 W=7.5e-07 $X=1360 $Y=345 $D=0
M2 7 A1 ZN VSS N L=1.8e-07 W=7.5e-07 $X=2080 $Y=345 $D=0
M3 VSS A2 7 VSS N L=1.8e-07 W=7.5e-07 $X=2690 $Y=345 $D=0
M4 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=740 $Y=2205 $D=16
M5 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1460 $Y=2205 $D=16
M6 ZN A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=2260 $Y=2205 $D=16
M7 VDD A2 ZN VDD P L=1.8e-07 W=6.85e-07 $X=2980 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IIND4D1BWP7T A1 B1 B2 ZN VSS VDD A2
** N=12 EP=7 IP=0 FDC=12
M0 8 A1 VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=345 $D=0
M1 10 8 ZN VSS N L=1.8e-07 W=1e-06 $X=2055 $Y=345 $D=0
M2 11 B1 10 VSS N L=1.8e-07 W=1e-06 $X=2665 $Y=345 $D=0
M3 12 B2 11 VSS N L=1.8e-07 W=1e-06 $X=3275 $Y=345 $D=0
M4 VSS 9 12 VSS N L=1.8e-07 W=1e-06 $X=3885 $Y=345 $D=0
M5 9 A2 VSS VSS N L=1.8e-07 W=5e-07 $X=4800 $Y=345 $D=0
M6 VDD A1 8 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2890 $D=16
M7 ZN 8 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M8 VDD B1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M9 ZN B2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3165 $Y=2205 $D=16
M10 VDD 9 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3885 $Y=2205 $D=16
M11 9 A2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=4800 $Y=2890 $D=16
.ENDS
***************************************
.SUBCKT INR2XD1BWP7T A1 ZN B1 VSS VDD
** N=7 EP=5 IP=0 FDC=8
M0 VSS A1 7 VSS N L=1.8e-07 W=1e-06 $X=640 $Y=345 $D=0
M1 ZN 7 VSS VSS N L=1.8e-07 W=1e-06 $X=1640 $Y=345 $D=0
M2 VSS B1 ZN VSS N L=1.8e-07 W=1e-06 $X=2535 $Y=345 $D=0
M3 VDD A1 7 VDD P L=1.8e-07 W=1.37e-06 $X=640 $Y=2205 $D=16
M4 6 7 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1520 $Y=2205 $D=16
M5 ZN B1 6 VDD P L=1.8e-07 W=1.37e-06 $X=2240 $Y=2205 $D=16
M6 6 B1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2960 $Y=2205 $D=16
M7 VDD 7 6 VDD P L=1.8e-07 W=1.37e-06 $X=3680 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INVD1P5BWP7T I ZN VSS VDD
** N=4 EP=4 IP=0 FDC=4
M0 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=670 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=5e-07 $X=1440 $Y=345 $D=0
M2 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=670 $Y=2205 $D=16
M3 VDD I ZN VDD P L=1.8e-07 W=6.85e-07 $X=1440 $Y=2890 $D=16
.ENDS
***************************************
.SUBCKT AOI211XD2BWP7T C VDD B A2 VSS ZN A1
** N=10 EP=7 IP=0 FDC=24
M0 ZN B VSS VSS N L=1.8e-07 W=1e-06 $X=720 $Y=345 $D=0
M1 VSS C ZN VSS N L=1.8e-07 W=1e-06 $X=2960 $Y=345 $D=0
M2 ZN C VSS VSS N L=1.8e-07 W=1e-06 $X=3760 $Y=345 $D=0
M3 VSS B ZN VSS N L=1.8e-07 W=1e-06 $X=4480 $Y=345 $D=0
M4 VSS A2 10 VSS N L=1.8e-07 W=1e-06 $X=8220 $Y=345 $D=0
M5 10 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=9020 $Y=345 $D=0
M6 ZN A1 10 VSS N L=1.8e-07 W=1e-06 $X=9800 $Y=345 $D=0
M7 10 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=10520 $Y=345 $D=0
M8 9 B 8 VDD P L=1.8e-07 W=1.37e-06 $X=720 $Y=2205 $D=16
M9 VDD C 9 VDD P L=1.8e-07 W=1.37e-06 $X=1440 $Y=2205 $D=16
M10 9 C VDD VDD P L=1.8e-07 W=1.37e-06 $X=2240 $Y=2205 $D=16
M11 VDD C 9 VDD P L=1.8e-07 W=1.37e-06 $X=2960 $Y=2205 $D=16
M12 9 C VDD VDD P L=1.8e-07 W=1.37e-06 $X=3760 $Y=2205 $D=16
M13 8 B 9 VDD P L=1.8e-07 W=1.37e-06 $X=4480 $Y=2205 $D=16
M14 9 B 8 VDD P L=1.8e-07 W=1.37e-06 $X=5200 $Y=2205 $D=16
M15 8 B 9 VDD P L=1.8e-07 W=1.37e-06 $X=5920 $Y=2205 $D=16
M16 ZN A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=6720 $Y=2205 $D=16
M17 8 A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=7480 $Y=2205 $D=16
M18 ZN A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=8240 $Y=2205 $D=16
M19 8 A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=9020 $Y=2205 $D=16
M20 ZN A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=9800 $Y=2205 $D=16
M21 8 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=10560 $Y=2205 $D=16
M22 ZN A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=11280 $Y=2205 $D=16
M23 8 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=12005 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR2XD2BWP7T A2 VDD VSS ZN A1
** N=6 EP=5 IP=0 FDC=12
M0 ZN A2 VSS VSS N L=1.8e-07 W=1e-06 $X=2100 $Y=345 $D=0
M1 VSS A2 ZN VSS N L=1.8e-07 W=1e-06 $X=2820 $Y=345 $D=0
M2 ZN A1 VSS VSS N L=1.8e-07 W=1e-06 $X=3540 $Y=345 $D=0
M3 VSS A1 ZN VSS N L=1.8e-07 W=1e-06 $X=4260 $Y=345 $D=0
M4 VDD A2 6 VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M5 6 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1380 $Y=2205 $D=16
M6 VDD A2 6 VDD P L=1.8e-07 W=1.37e-06 $X=2100 $Y=2205 $D=16
M7 6 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2820 $Y=2205 $D=16
M8 ZN A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=3540 $Y=2205 $D=16
M9 6 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4260 $Y=2205 $D=16
M10 ZN A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=4980 $Y=2205 $D=16
M11 6 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=5700 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_22 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480
+ 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500
+ 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520
+ 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540
+ 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560
+ 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580
+ 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600
+ 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620
+ 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640
+ 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660
+ 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680
+ 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698
** N=1183 EP=698 IP=6438 FDC=9254
M0 1181 959 1 1 N L=1.8e-07 W=1e-06 $X=180820 $Y=380985 $D=0
M1 979 939 1181 1 N L=1.8e-07 W=1e-06 $X=181540 $Y=380985 $D=0
M2 1 977 979 1 N L=1.8e-07 W=1e-06 $X=182380 $Y=380985 $D=0
M3 312 979 1 1 N L=1.8e-07 W=1e-06 $X=183220 $Y=380985 $D=0
M4 239 980 1 1 N L=1.8e-07 W=6.85e-07 $X=206740 $Y=388885 $D=0
M5 1 980 239 1 N L=1.8e-07 W=8.9e-07 $X=207460 $Y=388885 $D=0
M6 350 1012 1 1 N L=1.8e-07 W=1e-06 $X=208780 $Y=396665 $D=0
M7 1 1012 350 1 N L=1.8e-07 W=1e-06 $X=209515 $Y=396665 $D=0
M8 1008 962 1 1 N L=1.8e-07 W=1e-06 $X=210235 $Y=396665 $D=0
M9 1012 256 1008 1 N L=1.8e-07 W=1e-06 $X=210955 $Y=396665 $D=0
M10 1008 998 1012 1 N L=1.8e-07 W=1e-06 $X=211675 $Y=396665 $D=0
M11 1012 999 1008 1 N L=1.8e-07 W=1e-06 $X=212395 $Y=396665 $D=0
M12 979 959 974 2 P L=1.8e-07 W=1.37e-06 $X=180820 $Y=382845 $D=16
M13 974 939 979 2 P L=1.8e-07 W=1.37e-06 $X=181540 $Y=382845 $D=16
M14 2 977 974 2 P L=1.8e-07 W=1.37e-06 $X=182380 $Y=382845 $D=16
M15 312 979 2 2 P L=1.8e-07 W=1.37e-06 $X=183220 $Y=382845 $D=16
M16 2 980 239 2 P L=1.8e-07 W=1.37e-06 $X=206600 $Y=390685 $D=16
M17 239 980 2 2 P L=1.8e-07 W=1.37e-06 $X=207400 $Y=390685 $D=16
M18 2 980 239 2 P L=1.8e-07 W=1.37e-06 $X=208120 $Y=390685 $D=16
M19 350 1012 2 2 P L=1.8e-07 W=1.37e-06 $X=208780 $Y=398525 $D=16
M20 2 1012 350 2 P L=1.8e-07 W=1.37e-06 $X=209515 $Y=398525 $D=16
M21 1012 962 2 2 P L=1.8e-07 W=1.37e-06 $X=210280 $Y=398525 $D=16
M22 1182 256 1012 2 P L=1.8e-07 W=1.37e-06 $X=211055 $Y=398525 $D=16
M23 1183 998 1182 2 P L=1.8e-07 W=1.37e-06 $X=211710 $Y=398525 $D=16
M24 2 999 1183 2 P L=1.8e-07 W=1.37e-06 $X=212365 $Y=398525 $D=16
D25 1 980 DN AREA=2.037e-13 PJ=1.81e-06 $X=208720 $Y=389335 $D=32
X112 1 685 ANTENNABWP7T $T=471920 364960 0 180 $X=470510 $Y=360750
X113 1 686 ANTENNABWP7T $T=471920 372800 0 180 $X=470510 $Y=368590
X114 1 687 ANTENNABWP7T $T=471920 380640 0 180 $X=470510 $Y=376430
X115 1 690 ANTENNABWP7T $T=471920 388480 0 180 $X=470510 $Y=384270
X116 1 629 ANTENNABWP7T $T=471920 396320 0 180 $X=470510 $Y=392110
X117 1 630 ANTENNABWP7T $T=471920 404160 0 180 $X=470510 $Y=399950
X118 1 626 ANTENNABWP7T $T=471920 412000 0 180 $X=470510 $Y=407790
X119 1 628 ANTENNABWP7T $T=473040 364960 0 180 $X=471630 $Y=360750
X120 1 677 ANTENNABWP7T $T=473040 372800 0 180 $X=471630 $Y=368590
X121 1 663 ANTENNABWP7T $T=473040 380640 0 180 $X=471630 $Y=376430
X122 1 491 ANTENNABWP7T $T=473040 388480 0 180 $X=471630 $Y=384270
X123 1 693 ANTENNABWP7T $T=473040 396320 0 180 $X=471630 $Y=392110
X124 1 694 ANTENNABWP7T $T=473040 404160 0 180 $X=471630 $Y=399950
X125 1 418 ANTENNABWP7T $T=473040 412000 0 180 $X=471630 $Y=407790
X126 1 695 ANTENNABWP7T $T=473040 357120 0 0 $X=472750 $Y=356885
X127 1 510 ANTENNABWP7T $T=474160 364960 0 180 $X=472750 $Y=360750
X128 1 678 ANTENNABWP7T $T=473040 364960 0 0 $X=472750 $Y=364725
X129 1 676 ANTENNABWP7T $T=474160 372800 0 180 $X=472750 $Y=368590
X130 1 679 ANTENNABWP7T $T=473040 372800 0 0 $X=472750 $Y=372565
X131 1 548 ANTENNABWP7T $T=474160 380640 0 180 $X=472750 $Y=376430
X132 1 658 ANTENNABWP7T $T=474160 388480 0 180 $X=472750 $Y=384270
X133 1 644 ANTENNABWP7T $T=473040 388480 0 0 $X=472750 $Y=388245
X134 1 621 ANTENNABWP7T $T=474160 396320 0 180 $X=472750 $Y=392110
X135 1 697 ANTENNABWP7T $T=473040 396320 0 0 $X=472750 $Y=396085
X136 1 669 ANTENNABWP7T $T=474160 404160 0 180 $X=472750 $Y=399950
X137 1 573 ANTENNABWP7T $T=473040 404160 0 0 $X=472750 $Y=403925
X138 1 479 ANTENNABWP7T $T=474160 412000 0 180 $X=472750 $Y=407790
X139 1 698 ANTENNABWP7T $T=473040 412000 0 0 $X=472750 $Y=411765
X140 1 613 680 ICV_1 $T=469680 380640 0 0 $X=469390 $Y=380405
X141 1 683 692 ICV_1 $T=470800 357120 0 0 $X=470510 $Y=356885
X142 1 457 688 ICV_1 $T=470800 364960 0 0 $X=470510 $Y=364725
X143 1 665 689 ICV_1 $T=470800 372800 0 0 $X=470510 $Y=372565
X144 1 637 691 ICV_1 $T=470800 388480 0 0 $X=470510 $Y=388245
X145 1 642 560 ICV_1 $T=470800 396320 0 0 $X=470510 $Y=396085
X146 1 655 662 ICV_1 $T=470800 404160 0 0 $X=470510 $Y=403925
X147 1 684 506 ICV_1 $T=470800 412000 0 0 $X=470510 $Y=411765
X148 1 671 696 ICV_1 $T=471920 380640 0 0 $X=471630 $Y=380405
X228 795 1 2 16 CKBD1BWP7T $T=23920 396320 1 0 $X=23630 $Y=392110
X229 812 1 2 64 CKBD1BWP7T $T=46880 372800 1 0 $X=46590 $Y=368590
X230 265 1 2 942 CKBD1BWP7T $T=163920 364960 1 0 $X=163630 $Y=360750
X231 298 1 2 301 CKBD1BWP7T $T=176800 357120 0 0 $X=176510 $Y=356885
X232 1055 1 2 434 CKBD1BWP7T $T=278720 388480 1 180 $X=276190 $Y=388245
X233 1057 1 2 1056 CKBD1BWP7T $T=280400 372800 0 180 $X=277870 $Y=368590
X234 1108 1 2 1060 CKBD1BWP7T $T=353200 396320 1 0 $X=352910 $Y=392110
X235 548 1 2 545 CKBD1BWP7T $T=376160 372800 1 180 $X=373630 $Y=372565
X236 615 1 2 519 CKBD1BWP7T $T=434960 357120 1 180 $X=432430 $Y=356885
X237 550 1 2 618 CKBD1BWP7T $T=438880 388480 0 180 $X=436350 $Y=384270
X238 612 1 2 602 CKBD1BWP7T $T=442800 388480 0 180 $X=440270 $Y=384270
X239 629 1 2 625 CKBD1BWP7T $T=446720 388480 0 180 $X=444190 $Y=384270
X240 635 1 2 1170 CKBD1BWP7T $T=447840 380640 0 180 $X=445310 $Y=376430
X241 646 1 2 1150 CKBD1BWP7T $T=460720 357120 0 0 $X=460430 $Y=356885
X242 414 1 2 645 CKBD1BWP7T $T=462960 364960 0 180 $X=460430 $Y=360750
X243 647 1 2 1081 CKBD1BWP7T $T=463520 388480 0 180 $X=460990 $Y=384270
X244 663 1 2 660 CKBD1BWP7T $T=468560 380640 0 180 $X=466030 $Y=376430
X245 676 1 2 674 CKBD1BWP7T $T=470800 357120 1 180 $X=468270 $Y=356885
X246 681 1 2 580 CKBD1BWP7T $T=470800 388480 0 180 $X=468270 $Y=384270
X247 682 1 2 672 CKBD1BWP7T $T=470800 404160 0 180 $X=468270 $Y=399950
X248 788 1 2 801 INVD0BWP7T $T=23360 388480 1 0 $X=23070 $Y=384270
X249 45 1 2 52 INVD0BWP7T $T=41840 412000 0 0 $X=41550 $Y=411765
X250 70 1 2 827 INVD0BWP7T $T=50240 412000 1 0 $X=49950 $Y=407790
X251 833 1 2 87 INVD0BWP7T $T=58640 364960 0 180 $X=56670 $Y=360750
X252 817 1 2 108 INVD0BWP7T $T=62000 412000 1 0 $X=61710 $Y=407790
X253 26 1 2 105 INVD0BWP7T $T=64240 404160 0 180 $X=62270 $Y=399950
X254 93 1 2 111 INVD0BWP7T $T=65920 412000 1 180 $X=63950 $Y=411765
X255 39 1 2 846 INVD0BWP7T $T=67040 357120 0 0 $X=66750 $Y=356885
X256 158 1 2 155 INVD0BWP7T $T=87760 412000 0 180 $X=85790 $Y=407790
X257 862 1 2 856 INVD0BWP7T $T=90560 380640 1 180 $X=88590 $Y=380405
X258 186 1 2 875 INVD0BWP7T $T=102880 357120 0 0 $X=102590 $Y=356885
X259 20 1 2 885 INVD0BWP7T $T=109040 388480 0 180 $X=107070 $Y=384270
X260 871 1 2 887 INVD0BWP7T $T=123600 412000 0 180 $X=121630 $Y=407790
X261 187 1 2 898 INVD0BWP7T $T=129760 357120 1 180 $X=127790 $Y=356885
X262 900 1 2 911 INVD0BWP7T $T=137040 396320 1 0 $X=136750 $Y=392110
X263 236 1 2 914 INVD0BWP7T $T=147680 364960 0 180 $X=145710 $Y=360750
X264 231 1 2 941 INVD0BWP7T $T=163920 412000 1 0 $X=163630 $Y=407790
X265 922 1 2 946 INVD0BWP7T $T=165040 372800 1 0 $X=164750 $Y=368590
X266 279 1 2 274 INVD0BWP7T $T=169520 404160 0 180 $X=167550 $Y=399950
X267 968 1 2 295 INVD0BWP7T $T=176800 388480 0 180 $X=174830 $Y=384270
X268 306 1 2 938 INVD0BWP7T $T=180160 404160 1 180 $X=178190 $Y=403925
X269 313 1 2 299 INVD0BWP7T $T=183520 412000 1 0 $X=183230 $Y=407790
X270 963 1 2 987 INVD0BWP7T $T=188560 364960 0 0 $X=188270 $Y=364725
X271 989 1 2 330 INVD0BWP7T $T=191920 380640 1 180 $X=189950 $Y=380405
X272 991 1 2 989 INVD0BWP7T $T=192480 380640 0 180 $X=190510 $Y=376430
X273 1014 1 2 339 INVD0BWP7T $T=215440 364960 1 180 $X=213470 $Y=364725
X274 995 1 2 357 INVD0BWP7T $T=215440 396320 0 180 $X=213470 $Y=392110
X275 358 1 2 1019 INVD0BWP7T $T=223840 412000 1 0 $X=223550 $Y=407790
X276 1054 1 2 1042 INVD0BWP7T $T=272560 364960 0 180 $X=270590 $Y=360750
X277 446 1 2 1046 INVD0BWP7T $T=291600 364960 1 180 $X=289630 $Y=364725
X278 1067 1 2 1073 INVD0BWP7T $T=302240 396320 1 0 $X=301950 $Y=392110
X279 1082 1 2 1077 INVD0BWP7T $T=320160 380640 0 180 $X=318190 $Y=376430
X280 1090 1 2 1091 INVD0BWP7T $T=331920 388480 0 0 $X=331630 $Y=388245
X281 1079 1 2 1093 INVD0BWP7T $T=332480 404160 1 0 $X=332190 $Y=399950
X282 1097 1 2 1106 INVD0BWP7T $T=339760 372800 0 0 $X=339470 $Y=372565
X283 1101 1 2 1104 INVD0BWP7T $T=348160 396320 1 0 $X=347870 $Y=392110
X284 1113 1 2 1114 INVD0BWP7T $T=358240 396320 0 0 $X=357950 $Y=396085
X285 1081 1 2 1121 INVD0BWP7T $T=366640 396320 1 180 $X=364670 $Y=396085
X286 539 1 2 1127 INVD0BWP7T $T=377280 412000 1 0 $X=376990 $Y=407790
X287 571 1 2 1136 INVD0BWP7T $T=392400 372800 0 180 $X=390430 $Y=368590
X288 582 1 2 1145 INVD0BWP7T $T=398000 364960 1 0 $X=397710 $Y=360750
X289 1141 1 2 1154 INVD0BWP7T $T=406960 396320 0 0 $X=406670 $Y=396085
X290 633 1 2 622 INVD0BWP7T $T=446160 364960 0 180 $X=444190 $Y=360750
X291 641 1 2 1172 INVD0BWP7T $T=457920 404160 0 0 $X=457630 $Y=403925
X292 1150 1 2 656 INVD0BWP7T $T=462960 364960 1 0 $X=462670 $Y=360750
X293 653 1 2 666 INVD0BWP7T $T=466880 357120 0 0 $X=466590 $Y=356885
X294 643 1 2 1174 INVD0BWP7T $T=469680 396320 1 180 $X=467710 $Y=396085
X295 281 285 1 2 BUFFD1P5BWP7T $T=169520 357120 0 0 $X=169230 $Y=356885
X296 1031 400 1 2 BUFFD1P5BWP7T $T=239520 396320 0 180 $X=236430 $Y=392110
X297 1022 402 1 2 BUFFD1P5BWP7T $T=237840 380640 0 0 $X=237550 $Y=380405
X298 1061 441 1 2 BUFFD1P5BWP7T $T=282080 396320 0 180 $X=278990 $Y=392110
X299 1064 442 1 2 BUFFD1P5BWP7T $T=283200 412000 1 180 $X=280110 $Y=411765
X300 1066 445 1 2 BUFFD1P5BWP7T $T=294400 396320 0 180 $X=291310 $Y=392110
X301 1069 369 1 2 BUFFD1P5BWP7T $T=297200 404160 0 180 $X=294110 $Y=399950
X302 1124 549 1 2 BUFFD1P5BWP7T $T=378400 396320 0 180 $X=375310 $Y=392110
X303 630 623 1 2 BUFFD1P5BWP7T $T=446720 404160 0 180 $X=443630 $Y=399950
X304 637 634 1 2 BUFFD1P5BWP7T $T=449520 364960 0 180 $X=446430 $Y=360750
X305 642 638 1 2 BUFFD1P5BWP7T $T=460720 396320 0 180 $X=457630 $Y=392110
X306 644 639 1 2 BUFFD1P5BWP7T $T=461280 380640 1 180 $X=458190 $Y=380405
X307 658 652 1 2 BUFFD1P5BWP7T $T=466880 380640 1 180 $X=463790 $Y=380405
X308 665 657 1 2 BUFFD1P5BWP7T $T=468560 364960 1 180 $X=465470 $Y=364725
X309 671 661 1 2 BUFFD1P5BWP7T $T=469680 380640 1 180 $X=466590 $Y=380405
X310 677 659 1 2 BUFFD1P5BWP7T $T=470800 364960 0 180 $X=467710 $Y=360750
X311 679 667 1 2 BUFFD1P5BWP7T $T=470800 372800 0 180 $X=467710 $Y=368590
X312 1134 1 2 664 INVD3BWP7T $T=464640 396320 0 0 $X=464350 $Y=396085
X313 1175 1 2 675 INVD3BWP7T $T=466880 388480 0 0 $X=466590 $Y=388245
X314 416 418 2 1 418 1038 416 MAOI22D0BWP7T $T=260240 388480 0 0 $X=259950 $Y=388245
X315 462 458 2 1 462 1050 458 MAOI22D0BWP7T $T=302240 396320 0 180 $X=298030 $Y=392110
X316 450 479 2 1 479 1075 450 MAOI22D0BWP7T $T=314000 404160 0 180 $X=309790 $Y=399950
X317 460 506 2 1 506 1084 460 MAOI22D0BWP7T $T=324640 404160 1 180 $X=320430 $Y=403925
X318 514 510 2 1 514 1076 510 MAOI22D0BWP7T $T=338640 364960 1 180 $X=334430 $Y=364725
X382 474 540 474 540 1062 1 2 MAOI22D2BWP7T $T=363840 412000 0 180 $X=357390 $Y=407790
X383 880 1 2 197 BUFFD1BWP7T $T=106240 364960 0 0 $X=105950 $Y=364725
X384 917 1 2 926 BUFFD1BWP7T $T=144320 396320 0 0 $X=144030 $Y=396085
X385 924 1 2 919 BUFFD1BWP7T $T=146560 412000 1 180 $X=144030 $Y=411765
X386 272 1 2 950 BUFFD1BWP7T $T=165600 357120 0 0 $X=165310 $Y=356885
X387 1120 1 2 1118 BUFFD1BWP7T $T=366080 396320 0 180 $X=363550 $Y=392110
X388 605 1 2 603 BUFFD1BWP7T $T=425440 404160 1 180 $X=422910 $Y=403925
X389 607 1 2 1165 BUFFD1BWP7T $T=427120 364960 1 0 $X=426830 $Y=360750
X390 571 1 2 640 BUFFD1BWP7T $T=460720 357120 1 180 $X=458190 $Y=356885
X391 678 1 2 673 BUFFD1BWP7T $T=470800 364960 1 180 $X=468270 $Y=364725
X392 680 1 2 670 BUFFD1BWP7T $T=470800 380640 0 180 $X=468270 $Y=376430
X393 1 2 DCAP4BWP7T $T=21120 388480 1 0 $X=20830 $Y=384270
X394 1 2 DCAP4BWP7T $T=39600 396320 0 0 $X=39310 $Y=396085
X395 1 2 DCAP4BWP7T $T=58080 396320 0 0 $X=57790 $Y=396085
X396 1 2 DCAP4BWP7T $T=91680 404160 1 0 $X=91390 $Y=399950
X397 1 2 DCAP4BWP7T $T=99520 404160 1 0 $X=99230 $Y=399950
X398 1 2 DCAP4BWP7T $T=123600 380640 0 0 $X=123310 $Y=380405
X399 1 2 DCAP4BWP7T $T=134240 364960 0 0 $X=133950 $Y=364725
X400 1 2 DCAP4BWP7T $T=147120 372800 1 0 $X=146830 $Y=368590
X401 1 2 DCAP4BWP7T $T=157760 372800 1 0 $X=157470 $Y=368590
X402 1 2 DCAP4BWP7T $T=157760 412000 0 0 $X=157470 $Y=411765
X403 1 2 DCAP4BWP7T $T=182400 380640 1 0 $X=182110 $Y=376430
X404 1 2 DCAP4BWP7T $T=213200 380640 1 0 $X=212910 $Y=376430
X405 1 2 DCAP4BWP7T $T=232800 364960 0 0 $X=232510 $Y=364725
X406 1 2 DCAP4BWP7T $T=249600 364960 1 0 $X=249310 $Y=360750
X407 1 2 DCAP4BWP7T $T=249600 372800 1 0 $X=249310 $Y=368590
X408 1 2 DCAP4BWP7T $T=249600 380640 0 0 $X=249310 $Y=380405
X409 1 2 DCAP4BWP7T $T=249600 404160 1 0 $X=249310 $Y=399950
X410 1 2 DCAP4BWP7T $T=291600 412000 1 0 $X=291310 $Y=407790
X411 1 2 DCAP4BWP7T $T=307280 372800 1 0 $X=306990 $Y=368590
X412 1 2 DCAP4BWP7T $T=314000 388480 0 0 $X=313710 $Y=388245
X413 1 2 DCAP4BWP7T $T=325760 396320 0 0 $X=325470 $Y=396085
X414 1 2 DCAP4BWP7T $T=333600 357120 0 0 $X=333310 $Y=356885
X415 1 2 DCAP4BWP7T $T=333600 412000 1 0 $X=333310 $Y=407790
X416 1 2 DCAP4BWP7T $T=338080 412000 0 0 $X=337790 $Y=411765
X417 1 2 DCAP4BWP7T $T=352640 364960 1 0 $X=352350 $Y=360750
X418 1 2 DCAP4BWP7T $T=359360 404160 1 0 $X=359070 $Y=399950
X419 1 2 DCAP4BWP7T $T=367760 388480 1 0 $X=367470 $Y=384270
X420 1 2 DCAP4BWP7T $T=367760 388480 0 0 $X=367470 $Y=388245
X421 1 2 DCAP4BWP7T $T=375600 388480 0 0 $X=375310 $Y=388245
X422 1 2 DCAP4BWP7T $T=382880 396320 1 0 $X=382590 $Y=392110
X423 1 2 DCAP4BWP7T $T=394080 388480 0 0 $X=393790 $Y=388245
X424 1 2 DCAP4BWP7T $T=417600 388480 1 0 $X=417310 $Y=384270
X425 1 2 DCAP4BWP7T $T=428800 357120 0 0 $X=428510 $Y=356885
X426 1 2 DCAP4BWP7T $T=434960 357120 0 0 $X=434670 $Y=356885
X427 1 2 DCAP4BWP7T $T=435520 364960 0 0 $X=435230 $Y=364725
X428 1 2 DCAP4BWP7T $T=451760 380640 0 0 $X=451470 $Y=380405
X429 1 2 DCAP4BWP7T $T=455120 404160 1 0 $X=454830 $Y=399950
X430 1 2 DCAP4BWP7T $T=463520 364960 0 0 $X=463230 $Y=364725
X431 1 2 ICV_3 $T=25600 412000 1 0 $X=25310 $Y=407790
X432 1 2 ICV_3 $T=31200 357120 0 0 $X=30910 $Y=356885
X433 1 2 ICV_3 $T=31200 380640 1 0 $X=30910 $Y=376430
X434 1 2 ICV_3 $T=31200 396320 0 0 $X=30910 $Y=396085
X435 1 2 ICV_3 $T=31200 404160 1 0 $X=30910 $Y=399950
X436 1 2 ICV_3 $T=35120 412000 1 0 $X=34830 $Y=407790
X437 1 2 ICV_3 $T=39600 372800 1 0 $X=39310 $Y=368590
X438 1 2 ICV_3 $T=48000 412000 0 0 $X=47710 $Y=411765
X439 1 2 ICV_3 $T=52480 372800 1 0 $X=52190 $Y=368590
X440 1 2 ICV_3 $T=57520 372800 1 0 $X=57230 $Y=368590
X441 1 2 ICV_3 $T=73200 364960 0 0 $X=72910 $Y=364725
X442 1 2 ICV_3 $T=115200 372800 1 0 $X=114910 $Y=368590
X443 1 2 ICV_3 $T=115200 388480 1 0 $X=114910 $Y=384270
X444 1 2 ICV_3 $T=115200 404160 0 0 $X=114910 $Y=403925
X445 1 2 ICV_3 $T=115200 412000 1 0 $X=114910 $Y=407790
X446 1 2 ICV_3 $T=119120 364960 1 0 $X=118830 $Y=360750
X447 1 2 ICV_3 $T=119120 380640 1 0 $X=118830 $Y=376430
X448 1 2 ICV_3 $T=128640 412000 1 0 $X=128350 $Y=407790
X449 1 2 ICV_3 $T=148240 380640 1 0 $X=147950 $Y=376430
X450 1 2 ICV_3 $T=157200 357120 0 0 $X=156910 $Y=356885
X451 1 2 ICV_3 $T=157200 396320 1 0 $X=156910 $Y=392110
X452 1 2 ICV_3 $T=157200 396320 0 0 $X=156910 $Y=396085
X453 1 2 ICV_3 $T=161120 380640 1 0 $X=160830 $Y=376430
X454 1 2 ICV_3 $T=185760 364960 0 0 $X=185470 $Y=364725
X455 1 2 ICV_3 $T=199200 372800 1 0 $X=198910 $Y=368590
X456 1 2 ICV_3 $T=199200 380640 1 0 $X=198910 $Y=376430
X457 1 2 ICV_3 $T=199200 396320 1 0 $X=198910 $Y=392110
X458 1 2 ICV_3 $T=199200 396320 0 0 $X=198910 $Y=396085
X459 1 2 ICV_3 $T=227760 380640 0 0 $X=227470 $Y=380405
X460 1 2 ICV_3 $T=228880 404160 0 0 $X=228590 $Y=403925
X461 1 2 ICV_3 $T=258560 364960 0 0 $X=258270 $Y=364725
X462 1 2 ICV_3 $T=275360 372800 1 0 $X=275070 $Y=368590
X463 1 2 ICV_3 $T=283200 364960 0 0 $X=282910 $Y=364725
X464 1 2 ICV_3 $T=283200 412000 0 0 $X=282910 $Y=411765
X465 1 2 ICV_3 $T=291600 404160 1 0 $X=291310 $Y=399950
X466 1 2 ICV_3 $T=315680 380640 1 0 $X=315390 $Y=376430
X467 1 2 ICV_3 $T=325200 357120 0 0 $X=324910 $Y=356885
X468 1 2 ICV_3 $T=325200 364960 1 0 $X=324910 $Y=360750
X469 1 2 ICV_3 $T=329120 388480 0 0 $X=328830 $Y=388245
X470 1 2 ICV_3 $T=333600 396320 0 0 $X=333310 $Y=396085
X471 1 2 ICV_3 $T=347040 412000 1 0 $X=346750 $Y=407790
X472 1 2 ICV_3 $T=367200 412000 0 0 $X=366910 $Y=411765
X473 1 2 ICV_3 $T=375600 396320 0 0 $X=375310 $Y=396085
X474 1 2 ICV_3 $T=409200 357120 0 0 $X=408910 $Y=356885
X475 1 2 ICV_3 $T=417600 396320 1 0 $X=417310 $Y=392110
X476 1 2 ICV_3 $T=433840 388480 1 0 $X=433550 $Y=384270
X477 1 2 ICV_3 $T=461280 380640 0 0 $X=460990 $Y=380405
X478 1 2 DCAP8BWP7T $T=29520 372800 0 0 $X=29230 $Y=372565
X479 1 2 DCAP8BWP7T $T=97840 404160 0 0 $X=97550 $Y=403925
X480 1 2 DCAP8BWP7T $T=112960 412000 0 0 $X=112670 $Y=411765
X481 1 2 DCAP8BWP7T $T=113520 404160 1 0 $X=113230 $Y=399950
X482 1 2 DCAP8BWP7T $T=119120 396320 0 0 $X=118830 $Y=396085
X483 1 2 DCAP8BWP7T $T=132560 380640 0 0 $X=132270 $Y=380405
X484 1 2 DCAP8BWP7T $T=142080 364960 0 0 $X=141790 $Y=364725
X485 1 2 DCAP8BWP7T $T=143760 357120 0 0 $X=143470 $Y=356885
X486 1 2 DCAP8BWP7T $T=144320 388480 1 0 $X=144030 $Y=384270
X487 1 2 DCAP8BWP7T $T=153280 372800 1 0 $X=152990 $Y=368590
X488 1 2 DCAP8BWP7T $T=153280 412000 0 0 $X=152990 $Y=411765
X489 1 2 DCAP8BWP7T $T=155520 364960 0 0 $X=155230 $Y=364725
X490 1 2 DCAP8BWP7T $T=166160 364960 1 0 $X=165870 $Y=360750
X491 1 2 DCAP8BWP7T $T=172320 357120 0 0 $X=172030 $Y=356885
X492 1 2 DCAP8BWP7T $T=185760 380640 0 0 $X=185470 $Y=380405
X493 1 2 DCAP8BWP7T $T=197520 357120 0 0 $X=197230 $Y=356885
X494 1 2 DCAP8BWP7T $T=221040 364960 1 0 $X=220750 $Y=360750
X495 1 2 DCAP8BWP7T $T=221600 380640 1 0 $X=221310 $Y=376430
X496 1 2 DCAP8BWP7T $T=235600 380640 1 0 $X=235310 $Y=376430
X497 1 2 DCAP8BWP7T $T=238960 412000 1 0 $X=238670 $Y=407790
X498 1 2 DCAP8BWP7T $T=239520 388480 1 0 $X=239230 $Y=384270
X499 1 2 DCAP8BWP7T $T=239520 396320 1 0 $X=239230 $Y=392110
X500 1 2 DCAP8BWP7T $T=245120 372800 1 0 $X=244830 $Y=368590
X501 1 2 DCAP8BWP7T $T=245120 412000 1 0 $X=244830 $Y=407790
X502 1 2 DCAP8BWP7T $T=255760 388480 0 0 $X=255470 $Y=388245
X503 1 2 DCAP8BWP7T $T=256320 372800 1 0 $X=256030 $Y=368590
X504 1 2 DCAP8BWP7T $T=261360 404160 0 0 $X=261070 $Y=403925
X505 1 2 DCAP8BWP7T $T=264160 380640 0 0 $X=263870 $Y=380405
X506 1 2 DCAP8BWP7T $T=280960 396320 0 0 $X=280670 $Y=396085
X507 1 2 DCAP8BWP7T $T=281520 404160 0 0 $X=281230 $Y=403925
X508 1 2 DCAP8BWP7T $T=287120 396320 0 0 $X=286830 $Y=396085
X509 1 2 DCAP8BWP7T $T=297200 404160 1 0 $X=296910 $Y=399950
X510 1 2 DCAP8BWP7T $T=301120 364960 1 0 $X=300830 $Y=360750
X511 1 2 DCAP8BWP7T $T=302240 404160 0 0 $X=301950 $Y=403925
X512 1 2 DCAP8BWP7T $T=311760 380640 0 0 $X=311470 $Y=380405
X513 1 2 DCAP8BWP7T $T=317360 372800 0 0 $X=317070 $Y=372565
X514 1 2 DCAP8BWP7T $T=321280 396320 0 0 $X=320990 $Y=396085
X515 1 2 DCAP8BWP7T $T=322960 380640 1 0 $X=322670 $Y=376430
X516 1 2 DCAP8BWP7T $T=322960 388480 0 0 $X=322670 $Y=388245
X517 1 2 DCAP8BWP7T $T=333600 388480 0 0 $X=333310 $Y=388245
X518 1 2 DCAP8BWP7T $T=344800 372800 1 0 $X=344510 $Y=368590
X519 1 2 DCAP8BWP7T $T=353760 396320 0 0 $X=353470 $Y=396085
X520 1 2 DCAP8BWP7T $T=355440 412000 0 0 $X=355150 $Y=411765
X521 1 2 DCAP8BWP7T $T=361600 364960 1 0 $X=361310 $Y=360750
X522 1 2 DCAP8BWP7T $T=362160 372800 1 0 $X=361870 $Y=368590
X523 1 2 DCAP8BWP7T $T=378400 396320 1 0 $X=378110 $Y=392110
X524 1 2 DCAP8BWP7T $T=380080 404160 0 0 $X=379790 $Y=403925
X525 1 2 DCAP8BWP7T $T=388480 357120 0 0 $X=388190 $Y=356885
X526 1 2 DCAP8BWP7T $T=393520 380640 1 0 $X=393230 $Y=376430
X527 1 2 DCAP8BWP7T $T=396880 404160 0 0 $X=396590 $Y=403925
X528 1 2 DCAP8BWP7T $T=404160 380640 0 0 $X=403870 $Y=380405
X529 1 2 DCAP8BWP7T $T=431040 396320 1 0 $X=430750 $Y=392110
X530 1 2 DCAP8BWP7T $T=447280 380640 0 0 $X=446990 $Y=380405
X531 1 2 DCAP8BWP7T $T=448960 372800 1 0 $X=448670 $Y=368590
X532 1 2 DCAP8BWP7T $T=449520 364960 1 0 $X=449230 $Y=360750
X533 1 2 DCAP8BWP7T $T=449520 372800 0 0 $X=449230 $Y=372565
X534 2 1 DCAPBWP7T $T=21120 372800 1 0 $X=20830 $Y=368590
X535 2 1 DCAPBWP7T $T=21120 380640 1 0 $X=20830 $Y=376430
X536 2 1 DCAPBWP7T $T=32320 404160 0 0 $X=32030 $Y=403925
X537 2 1 DCAPBWP7T $T=48560 412000 1 0 $X=48270 $Y=407790
X538 2 1 DCAPBWP7T $T=51920 412000 1 0 $X=51630 $Y=407790
X539 2 1 DCAPBWP7T $T=53600 404160 0 0 $X=53310 $Y=403925
X540 2 1 DCAPBWP7T $T=58640 364960 1 0 $X=58350 $Y=360750
X541 2 1 DCAPBWP7T $T=65920 412000 0 0 $X=65630 $Y=411765
X542 2 1 DCAPBWP7T $T=104000 372800 0 0 $X=103710 $Y=372565
X543 2 1 DCAPBWP7T $T=116320 396320 1 0 $X=116030 $Y=392110
X544 2 1 DCAPBWP7T $T=140400 388480 1 0 $X=140110 $Y=384270
X545 2 1 DCAPBWP7T $T=144320 380640 0 0 $X=144030 $Y=380405
X546 2 1 DCAPBWP7T $T=163360 404160 0 0 $X=163070 $Y=403925
X547 2 1 DCAPBWP7T $T=167840 357120 0 0 $X=167550 $Y=356885
X548 2 1 DCAPBWP7T $T=190240 404160 1 0 $X=189950 $Y=399950
X549 2 1 DCAPBWP7T $T=207600 388480 1 0 $X=207310 $Y=384270
X550 2 1 DCAPBWP7T $T=223280 412000 0 0 $X=222990 $Y=411765
X551 2 1 DCAPBWP7T $T=223840 388480 0 0 $X=223550 $Y=388245
X552 2 1 DCAPBWP7T $T=236160 380640 0 0 $X=235870 $Y=380405
X553 2 1 DCAPBWP7T $T=242320 412000 0 0 $X=242030 $Y=411765
X554 2 1 DCAPBWP7T $T=284320 357120 0 0 $X=284030 $Y=356885
X555 2 1 DCAPBWP7T $T=326320 388480 1 0 $X=326030 $Y=384270
X556 2 1 DCAPBWP7T $T=326320 404160 1 0 $X=326030 $Y=399950
X557 2 1 DCAPBWP7T $T=333600 380640 0 0 $X=333310 $Y=380405
X558 2 1 DCAPBWP7T $T=343680 412000 1 0 $X=343390 $Y=407790
X559 2 1 DCAPBWP7T $T=356000 412000 1 0 $X=355710 $Y=407790
X560 2 1 DCAPBWP7T $T=357680 380640 1 0 $X=357390 $Y=376430
X561 2 1 DCAPBWP7T $T=404160 357120 0 0 $X=403870 $Y=356885
X562 2 1 DCAPBWP7T $T=410320 364960 0 0 $X=410030 $Y=364725
X563 2 1 DCAPBWP7T $T=410320 388480 1 0 $X=410030 $Y=384270
X564 2 1 DCAPBWP7T $T=410320 404160 1 0 $X=410030 $Y=399950
X565 2 1 DCAPBWP7T $T=422080 380640 1 0 $X=421790 $Y=376430
X566 2 1 DCAPBWP7T $T=438880 388480 1 0 $X=438590 $Y=384270
X567 2 1 DCAPBWP7T $T=442800 388480 1 0 $X=442510 $Y=384270
X568 2 1 DCAPBWP7T $T=459600 388480 1 0 $X=459310 $Y=384270
X569 2 1 DCAPBWP7T $T=469120 412000 1 0 $X=468830 $Y=407790
X570 405 407 392 412 414 404 1 2 1032 AO222D0BWP7T $T=252400 364960 0 0 $X=252110 $Y=364725
X571 462 404 470 464 386 466 1 2 1037 AO222D0BWP7T $T=306720 372800 1 180 $X=300270 $Y=372565
X572 474 404 473 464 410 466 1 2 1041 AO222D0BWP7T $T=307840 404160 0 180 $X=301390 $Y=399950
X573 451 404 475 464 472 466 1 2 1033 AO222D0BWP7T $T=309520 380640 0 180 $X=303070 $Y=376430
X574 465 404 480 464 477 466 1 2 1034 AO222D0BWP7T $T=313440 396320 1 180 $X=306990 $Y=396085
X575 448 404 488 464 482 466 1 2 1043 AO222D0BWP7T $T=315680 380640 0 180 $X=309230 $Y=376430
X576 1081 404 491 464 486 466 1 2 1071 AO222D0BWP7T $T=317360 388480 0 180 $X=310910 $Y=384270
X577 405 518 412 1100 516 404 1 2 1102 AO222D0BWP7T $T=337520 364960 1 0 $X=337230 $Y=360750
X578 518 405 531 1100 536 404 1 2 537 AO222D0BWP7T $T=354320 357120 0 0 $X=354030 $Y=356885
X579 555 558 560 464 564 466 1 2 1135 AO222D0BWP7T $T=378400 396320 0 0 $X=378110 $Y=396085
X580 568 558 573 464 575 466 1 2 1139 AO222D0BWP7T $T=386800 396320 1 0 $X=386510 $Y=392110
X581 596 616 613 464 611 466 1 2 1164 AO222D0BWP7T $T=435520 364960 1 180 $X=429070 $Y=364725
X582 539 558 621 464 620 466 1 2 1167 AO222D0BWP7T $T=444480 396320 0 180 $X=438030 $Y=392110
X583 529 558 655 464 650 466 1 2 600 AO222D0BWP7T $T=467440 412000 1 180 $X=460990 $Y=411765
X584 643 558 662 464 654 466 1 2 649 AO222D0BWP7T $T=469120 412000 0 180 $X=462670 $Y=407790
X585 672 558 669 464 653 466 1 2 1171 AO222D0BWP7T $T=470800 404160 1 180 $X=464350 $Y=403925
X586 1 2 ICV_4 $T=21120 364960 0 0 $X=20830 $Y=364725
X587 1 2 ICV_4 $T=35120 380640 0 0 $X=34830 $Y=380405
X588 1 2 ICV_4 $T=39600 380640 1 0 $X=39310 $Y=376430
X589 1 2 ICV_4 $T=53600 404160 1 0 $X=53310 $Y=399950
X590 1 2 ICV_4 $T=119120 388480 1 0 $X=118830 $Y=384270
X591 1 2 ICV_4 $T=130320 372800 0 0 $X=130030 $Y=372565
X592 1 2 ICV_4 $T=130880 396320 0 0 $X=130590 $Y=396085
X593 1 2 ICV_4 $T=137040 412000 0 0 $X=136750 $Y=411765
X594 1 2 ICV_4 $T=148800 372800 0 0 $X=148510 $Y=372565
X595 1 2 ICV_4 $T=161120 372800 1 0 $X=160830 $Y=368590
X596 1 2 ICV_4 $T=161120 396320 1 0 $X=160830 $Y=392110
X597 1 2 ICV_4 $T=171200 388480 0 0 $X=170910 $Y=388245
X598 1 2 ICV_4 $T=221040 396320 0 0 $X=220750 $Y=396085
X599 1 2 ICV_4 $T=228880 372800 0 0 $X=228590 $Y=372565
X600 1 2 ICV_4 $T=228880 388480 1 0 $X=228590 $Y=384270
X601 1 2 ICV_4 $T=230000 412000 0 0 $X=229710 $Y=411765
X602 1 2 ICV_4 $T=240080 380640 1 0 $X=239790 $Y=376430
X603 1 2 ICV_4 $T=245120 388480 1 0 $X=244830 $Y=384270
X604 1 2 ICV_4 $T=245120 404160 0 0 $X=244830 $Y=403925
X605 1 2 ICV_4 $T=282080 396320 1 0 $X=281790 $Y=392110
X606 1 2 ICV_4 $T=282080 412000 1 0 $X=281790 $Y=407790
X607 1 2 ICV_4 $T=287120 372800 0 0 $X=286830 $Y=372565
X608 1 2 ICV_4 $T=287120 380640 1 0 $X=286830 $Y=376430
X609 1 2 ICV_4 $T=294400 396320 1 0 $X=294110 $Y=392110
X610 1 2 ICV_4 $T=305600 364960 1 0 $X=305310 $Y=360750
X611 1 2 ICV_4 $T=324080 412000 0 0 $X=323790 $Y=411765
X612 1 2 ICV_4 $T=333600 364960 1 0 $X=333310 $Y=360750
X613 1 2 ICV_4 $T=366080 396320 1 0 $X=365790 $Y=392110
X614 1 2 ICV_4 $T=371120 404160 1 0 $X=370830 $Y=399950
X615 1 2 ICV_4 $T=382320 364960 0 0 $X=382030 $Y=364725
X616 1 2 ICV_4 $T=392960 357120 0 0 $X=392670 $Y=356885
X617 1 2 ICV_4 $T=450080 364960 0 0 $X=449790 $Y=364725
X618 1 2 ICV_4 $T=450080 396320 0 0 $X=449790 $Y=396085
X619 372 1033 380 2 1 368 DFCNQD1BWP7T $T=260800 380640 0 180 $X=248190 $Y=376430
X620 372 1034 380 2 1 1029 DFCNQD1BWP7T $T=261360 388480 0 180 $X=248750 $Y=384270
X621 372 1035 380 2 1 1028 DFCNQD1BWP7T $T=261360 404160 1 180 $X=248750 $Y=403925
X622 372 415 380 2 1 1031 DFCNQD1BWP7T $T=262480 396320 1 180 $X=249870 $Y=396085
X623 372 1037 380 2 1 1030 DFCNQD1BWP7T $T=264160 380640 1 180 $X=251550 $Y=380405
X624 372 1039 380 2 1 1027 DFCNQD1BWP7T $T=265840 404160 0 180 $X=253230 $Y=399950
X625 372 1041 380 2 1 1026 DFCNQD1BWP7T $T=266400 396320 0 180 $X=253790 $Y=392110
X626 372 1043 380 2 1 413 DFCNQD1BWP7T $T=267520 372800 1 180 $X=254910 $Y=372565
X627 436 1045 380 2 1 1025 DFCNQD1BWP7T $T=278720 396320 0 180 $X=266110 $Y=392110
X628 436 1053 380 2 1 1036 DFCNQD1BWP7T $T=278720 404160 0 180 $X=266110 $Y=399950
X629 436 438 380 2 1 426 DFCNQD1BWP7T $T=280960 396320 1 180 $X=268350 $Y=396085
X630 436 1058 380 2 1 427 DFCNQD1BWP7T $T=281520 404160 1 180 $X=268910 $Y=403925
X631 436 459 380 2 1 1047 DFCNQD1BWP7T $T=302240 404160 1 180 $X=289630 $Y=403925
X632 436 463 380 2 1 1061 DFCNQD1BWP7T $T=303920 396320 1 180 $X=291310 $Y=396085
X633 436 467 380 2 1 449 DFCNQD1BWP7T $T=304480 412000 1 180 $X=291870 $Y=411765
X634 436 1071 380 2 1 1066 DFCNQD1BWP7T $T=305040 388480 1 180 $X=292430 $Y=388245
X635 436 468 380 2 1 1064 DFCNQD1BWP7T $T=306160 412000 0 180 $X=293550 $Y=407790
X636 436 499 380 2 1 1069 DFCNQD1BWP7T $T=321840 412000 0 180 $X=309230 $Y=407790
X637 436 504 494 2 1 484 DFCNQD1BWP7T $T=324080 412000 1 180 $X=311470 $Y=411765
X638 436 1135 532 2 1 1124 DFCNQD1BWP7T $T=387360 404160 0 180 $X=374750 $Y=399950
X639 436 1139 494 2 1 561 DFCNQD1BWP7T $T=396880 404160 1 180 $X=384270 $Y=403925
X640 436 1164 532 2 1 597 DFCNQD1BWP7T $T=432160 412000 0 180 $X=419550 $Y=407790
X641 436 1167 532 2 1 570 DFCNQD1BWP7T $T=435520 412000 1 180 $X=422910 $Y=411765
X642 436 614 532 2 1 604 DFCNQD1BWP7T $T=436080 380640 0 180 $X=423470 $Y=376430
X643 436 1171 532 2 1 1168 DFCNQD1BWP7T $T=448400 404160 1 180 $X=435790 $Y=403925
X644 436 636 532 2 1 619 DFCNQD1BWP7T $T=450080 364960 1 180 $X=437470 $Y=364725
X645 436 668 532 2 1 1173 DFCNQD1BWP7T $T=470800 372800 1 180 $X=458190 $Y=372565
X928 1 2 ICV_8 $T=20000 396320 1 0 $X=19710 $Y=392110
X929 1 2 ICV_8 $T=34000 357120 0 0 $X=33710 $Y=356885
X930 1 2 ICV_8 $T=34000 372800 0 0 $X=33710 $Y=372565
X931 1 2 ICV_8 $T=34000 388480 1 0 $X=33710 $Y=384270
X932 1 2 ICV_8 $T=34000 388480 0 0 $X=33710 $Y=388245
X933 1 2 ICV_8 $T=118000 404160 1 0 $X=117710 $Y=399950
X934 1 2 ICV_8 $T=118000 412000 1 0 $X=117710 $Y=407790
X935 1 2 ICV_8 $T=160000 357120 0 0 $X=159710 $Y=356885
X936 1 2 ICV_8 $T=160000 364960 1 0 $X=159710 $Y=360750
X937 1 2 ICV_8 $T=160000 404160 1 0 $X=159710 $Y=399950
X938 1 2 ICV_8 $T=160000 412000 0 0 $X=159710 $Y=411765
X939 1 2 ICV_8 $T=202000 380640 1 0 $X=201710 $Y=376430
X940 1 2 ICV_8 $T=202000 396320 1 0 $X=201710 $Y=392110
X941 1 2 ICV_8 $T=202000 396320 0 0 $X=201710 $Y=396085
X942 1 2 ICV_8 $T=286000 357120 0 0 $X=285710 $Y=356885
X943 1 2 ICV_8 $T=286000 364960 0 0 $X=285710 $Y=364725
X944 1 2 ICV_8 $T=286000 404160 0 0 $X=285710 $Y=403925
X945 1 2 ICV_8 $T=370000 364960 0 0 $X=369710 $Y=364725
X946 1 2 ICV_8 $T=412000 357120 0 0 $X=411710 $Y=356885
X947 1 2 ICV_8 $T=454000 404160 0 0 $X=453710 $Y=403925
X948 1 2 ICV_9 $T=20000 404160 1 0 $X=19710 $Y=399950
X949 1 2 ICV_9 $T=20000 412000 1 0 $X=19710 $Y=407790
X950 1 2 ICV_9 $T=34000 372800 1 0 $X=33710 $Y=368590
X951 1 2 ICV_9 $T=34000 380640 1 0 $X=33710 $Y=376430
X952 1 2 ICV_9 $T=34000 396320 1 0 $X=33710 $Y=392110
X953 1 2 ICV_9 $T=34000 396320 0 0 $X=33710 $Y=396085
X954 1 2 ICV_9 $T=34000 404160 1 0 $X=33710 $Y=399950
X955 1 2 ICV_9 $T=34000 404160 0 0 $X=33710 $Y=403925
X956 1 2 ICV_9 $T=118000 404160 0 0 $X=117710 $Y=403925
X957 1 2 ICV_9 $T=160000 364960 0 0 $X=159710 $Y=364725
X958 1 2 ICV_9 $T=202000 357120 0 0 $X=201710 $Y=356885
X959 1 2 ICV_9 $T=202000 372800 1 0 $X=201710 $Y=368590
X960 1 2 ICV_9 $T=202000 388480 1 0 $X=201710 $Y=384270
X961 1 2 ICV_9 $T=244000 357120 0 0 $X=243710 $Y=356885
X962 1 2 ICV_9 $T=244000 364960 1 0 $X=243710 $Y=360750
X963 1 2 ICV_9 $T=244000 364960 0 0 $X=243710 $Y=364725
X964 1 2 ICV_9 $T=244000 380640 0 0 $X=243710 $Y=380405
X965 1 2 ICV_9 $T=244000 388480 0 0 $X=243710 $Y=388245
X966 1 2 ICV_9 $T=244000 404160 1 0 $X=243710 $Y=399950
X967 1 2 ICV_9 $T=286000 388480 0 0 $X=285710 $Y=388245
X968 1 2 ICV_9 $T=286000 396320 1 0 $X=285710 $Y=392110
X969 1 2 ICV_9 $T=286000 404160 1 0 $X=285710 $Y=399950
X970 1 2 ICV_9 $T=286000 412000 1 0 $X=285710 $Y=407790
X971 1 2 ICV_9 $T=286000 412000 0 0 $X=285710 $Y=411765
X972 1 2 ICV_9 $T=328000 357120 0 0 $X=327710 $Y=356885
X973 1 2 ICV_9 $T=328000 364960 1 0 $X=327710 $Y=360750
X974 1 2 ICV_9 $T=328000 364960 0 0 $X=327710 $Y=364725
X975 1 2 ICV_9 $T=328000 372800 0 0 $X=327710 $Y=372565
X976 1 2 ICV_9 $T=328000 380640 0 0 $X=327710 $Y=380405
X977 1 2 ICV_9 $T=328000 388480 1 0 $X=327710 $Y=384270
X978 1 2 ICV_9 $T=328000 396320 1 0 $X=327710 $Y=392110
X979 1 2 ICV_9 $T=328000 396320 0 0 $X=327710 $Y=396085
X980 1 2 ICV_9 $T=328000 404160 0 0 $X=327710 $Y=403925
X981 1 2 ICV_9 $T=328000 412000 1 0 $X=327710 $Y=407790
X982 1 2 ICV_9 $T=370000 372800 1 0 $X=369710 $Y=368590
X983 1 2 ICV_9 $T=370000 388480 1 0 $X=369710 $Y=384270
X984 1 2 ICV_9 $T=370000 388480 0 0 $X=369710 $Y=388245
X985 1 2 ICV_9 $T=370000 396320 1 0 $X=369710 $Y=392110
X986 1 2 ICV_9 $T=370000 396320 0 0 $X=369710 $Y=396085
X987 1 2 ICV_9 $T=370000 412000 1 0 $X=369710 $Y=407790
X988 1 2 ICV_9 $T=370000 412000 0 0 $X=369710 $Y=411765
X989 1 2 ICV_9 $T=412000 364960 0 0 $X=411710 $Y=364725
X990 1 2 ICV_9 $T=412000 380640 0 0 $X=411710 $Y=380405
X991 1 2 ICV_9 $T=412000 388480 1 0 $X=411710 $Y=384270
X992 1 2 ICV_9 $T=412000 396320 1 0 $X=411710 $Y=392110
X993 1 2 ICV_9 $T=412000 404160 1 0 $X=411710 $Y=399950
X994 1 2 ICV_9 $T=412000 412000 1 0 $X=411710 $Y=407790
X995 1 2 ICV_9 $T=454000 364960 1 0 $X=453710 $Y=360750
X996 1 2 ICV_9 $T=454000 388480 1 0 $X=453710 $Y=384270
X997 1 2 ICV_9 $T=454000 388480 0 0 $X=453710 $Y=388245
X998 1 2 ICV_9 $T=454000 412000 1 0 $X=453710 $Y=407790
X1037 1 2 ICV_13 $T=21120 380640 0 0 $X=20830 $Y=380405
X1038 1 2 ICV_13 $T=30640 364960 0 0 $X=30350 $Y=364725
X1039 1 2 ICV_13 $T=30640 396320 1 0 $X=30350 $Y=392110
X1040 1 2 ICV_13 $T=35120 364960 1 0 $X=34830 $Y=360750
X1041 1 2 ICV_13 $T=35120 364960 0 0 $X=34830 $Y=364725
X1042 1 2 ICV_13 $T=97280 388480 0 0 $X=96990 $Y=388245
X1043 1 2 ICV_13 $T=119120 372800 1 0 $X=118830 $Y=368590
X1044 1 2 ICV_13 $T=119120 396320 1 0 $X=118830 $Y=392110
X1045 1 2 ICV_13 $T=123600 396320 0 0 $X=123310 $Y=396085
X1046 1 2 ICV_13 $T=123600 404160 0 0 $X=123310 $Y=403925
X1047 1 2 ICV_13 $T=138160 357120 0 0 $X=137870 $Y=356885
X1048 1 2 ICV_13 $T=146560 412000 0 0 $X=146270 $Y=411765
X1049 1 2 ICV_13 $T=149360 412000 1 0 $X=149070 $Y=407790
X1050 1 2 ICV_13 $T=156640 404160 1 0 $X=156350 $Y=399950
X1051 1 2 ICV_13 $T=156640 412000 1 0 $X=156350 $Y=407790
X1052 1 2 ICV_13 $T=161120 388480 1 0 $X=160830 $Y=384270
X1053 1 2 ICV_13 $T=161120 388480 0 0 $X=160830 $Y=388245
X1054 1 2 ICV_13 $T=161120 396320 0 0 $X=160830 $Y=396085
X1055 1 2 ICV_13 $T=170640 364960 1 0 $X=170350 $Y=360750
X1056 1 2 ICV_13 $T=198640 388480 1 0 $X=198350 $Y=384270
X1057 1 2 ICV_13 $T=203120 380640 0 0 $X=202830 $Y=380405
X1058 1 2 ICV_13 $T=203120 412000 1 0 $X=202830 $Y=407790
X1059 1 2 ICV_13 $T=203120 412000 0 0 $X=202830 $Y=411765
X1060 1 2 ICV_13 $T=212080 412000 0 0 $X=211790 $Y=411765
X1061 1 2 ICV_13 $T=225520 364960 1 0 $X=225230 $Y=360750
X1062 1 2 ICV_13 $T=226080 380640 1 0 $X=225790 $Y=376430
X1063 1 2 ICV_13 $T=240640 380640 0 0 $X=240350 $Y=380405
X1064 1 2 ICV_13 $T=240640 388480 0 0 $X=240350 $Y=388245
X1065 1 2 ICV_13 $T=245120 380640 1 0 $X=244830 $Y=376430
X1066 1 2 ICV_13 $T=249600 357120 0 0 $X=249310 $Y=356885
X1067 1 2 ICV_13 $T=260800 372800 1 0 $X=260510 $Y=368590
X1068 1 2 ICV_13 $T=264160 388480 0 0 $X=263870 $Y=388245
X1069 1 2 ICV_13 $T=265840 404160 0 0 $X=265550 $Y=403925
X1070 1 2 ICV_13 $T=282640 380640 1 0 $X=282350 $Y=376430
X1071 1 2 ICV_13 $T=303920 396320 0 0 $X=303630 $Y=396085
X1072 1 2 ICV_13 $T=308400 396320 1 0 $X=308110 $Y=392110
X1073 1 2 ICV_13 $T=314560 372800 1 0 $X=314270 $Y=368590
X1074 1 2 ICV_13 $T=329120 404160 1 0 $X=328830 $Y=399950
X1075 1 2 ICV_13 $T=338640 404160 1 0 $X=338350 $Y=399950
X1076 1 2 ICV_13 $T=342560 380640 1 0 $X=342270 $Y=376430
X1077 1 2 ICV_13 $T=347600 396320 0 0 $X=347310 $Y=396085
X1078 1 2 ICV_13 $T=349840 396320 1 0 $X=349550 $Y=392110
X1079 1 2 ICV_13 $T=366640 372800 1 0 $X=366350 $Y=368590
X1080 1 2 ICV_13 $T=366640 396320 0 0 $X=366350 $Y=396085
X1081 1 2 ICV_13 $T=377280 380640 1 0 $X=376990 $Y=376430
X1082 1 2 ICV_13 $T=392400 388480 1 0 $X=392110 $Y=384270
X1083 1 2 ICV_13 $T=408640 364960 1 0 $X=408350 $Y=360750
X1084 1 2 ICV_13 $T=408640 380640 0 0 $X=408350 $Y=380405
X1085 1 2 ICV_13 $T=408640 396320 0 0 $X=408350 $Y=396085
X1086 1 2 ICV_13 $T=413120 372800 1 0 $X=412830 $Y=368590
X1087 1 2 ICV_13 $T=417600 404160 1 0 $X=417310 $Y=399950
X1088 1 2 ICV_13 $T=427120 380640 0 0 $X=426830 $Y=380405
X1089 1 2 ICV_13 $T=432160 412000 1 0 $X=431870 $Y=407790
X1090 1 2 ICV_13 $T=455120 357120 0 0 $X=454830 $Y=356885
X1091 1 2 ICV_13 $T=455120 372800 0 0 $X=454830 $Y=372565
X1092 1 2 ICV_13 $T=459600 412000 1 0 $X=459310 $Y=407790
X1093 1 2 ICV_13 $T=463520 388480 0 0 $X=463230 $Y=388245
X1094 1 2 ICV_13 $T=464640 372800 1 0 $X=464350 $Y=368590
X1095 1 2 ICV_13 $T=467440 412000 0 0 $X=467150 $Y=411765
X1096 453 457 2 457 454 453 1 MAOI22D1BWP7T $T=301120 364960 0 180 $X=296350 $Y=360750
X1097 1136 574 2 574 1132 1136 1 MAOI22D1BWP7T $T=392400 364960 0 180 $X=387630 $Y=360750
X1098 622 628 2 628 1157 622 1 MAOI22D1BWP7T $T=448400 357120 1 180 $X=443630 $Y=356885
X1099 632 626 2 632 1153 626 1 MAOI22D1BWP7T $T=448960 412000 1 180 $X=444190 $Y=411765
X1100 1050 404 1 1039 423 2 IOA21D0BWP7T $T=270880 388480 1 180 $X=267230 $Y=388245
X1101 1062 404 1 1053 439 2 IOA21D0BWP7T $T=282080 412000 0 180 $X=278430 $Y=407790
X1102 483 404 1 1058 476 2 IOA21D0BWP7T $T=312320 404160 1 180 $X=308670 $Y=403925
X1103 14 1 2 799 INVD1BWP7T $T=25040 372800 1 0 $X=24750 $Y=368590
X1104 19 1 2 24 INVD1BWP7T $T=27280 357120 0 0 $X=26990 $Y=356885
X1105 35 1 2 46 INVD1BWP7T $T=43520 412000 0 180 $X=41550 $Y=407790
X1106 53 1 2 815 INVD1BWP7T $T=43520 412000 0 0 $X=43230 $Y=411765
X1107 807 1 2 61 INVD1BWP7T $T=45760 357120 0 0 $X=45470 $Y=356885
X1108 72 1 2 38 INVD1BWP7T $T=51920 357120 1 180 $X=49950 $Y=356885
X1109 802 1 2 103 INVD1BWP7T $T=62560 380640 0 180 $X=60590 $Y=376430
X1110 792 1 2 107 INVD1BWP7T $T=62000 388480 1 0 $X=61710 $Y=384270
X1111 127 1 2 824 INVD1BWP7T $T=71520 380640 0 0 $X=71230 $Y=380405
X1112 800 1 2 143 INVD1BWP7T $T=71520 412000 0 0 $X=71230 $Y=411765
X1113 150 1 2 145 INVD1BWP7T $T=85520 404160 0 180 $X=83550 $Y=399950
X1114 874 1 2 168 INVD1BWP7T $T=93360 364960 0 180 $X=91390 $Y=360750
X1115 814 1 2 834 INVD1BWP7T $T=91680 396320 0 0 $X=91390 $Y=396085
X1116 865 1 2 819 INVD1BWP7T $T=93360 396320 0 0 $X=93070 $Y=396085
X1117 861 1 2 178 INVD1BWP7T $T=99520 404160 0 180 $X=97550 $Y=399950
X1118 882 1 2 124 INVD1BWP7T $T=106800 372800 1 0 $X=106510 $Y=368590
X1119 199 1 2 42 INVD1BWP7T $T=110160 380640 0 180 $X=108190 $Y=376430
X1120 809 1 2 899 INVD1BWP7T $T=121920 364960 0 0 $X=121630 $Y=364725
X1121 904 1 2 889 INVD1BWP7T $T=130320 388480 0 180 $X=128350 $Y=384270
X1122 883 1 2 907 INVD1BWP7T $T=131440 404160 0 180 $X=129470 $Y=399950
X1123 884 1 2 849 INVD1BWP7T $T=138160 380640 0 180 $X=136190 $Y=376430
X1124 918 1 2 843 INVD1BWP7T $T=143200 380640 0 180 $X=141230 $Y=376430
X1125 935 1 2 934 INVD1BWP7T $T=155520 396320 0 0 $X=155230 $Y=396085
X1126 259 1 2 246 INVD1BWP7T $T=165600 357120 1 180 $X=163630 $Y=356885
X1127 269 1 2 260 INVD1BWP7T $T=165600 404160 0 180 $X=163630 $Y=399950
X1128 954 1 2 929 INVD1BWP7T $T=173440 380640 0 0 $X=173150 $Y=380405
X1129 945 1 2 287 INVD1BWP7T $T=175120 412000 0 180 $X=173150 $Y=407790
X1130 293 1 2 967 INVD1BWP7T $T=177920 404160 1 0 $X=177630 $Y=399950
X1131 305 1 2 270 INVD1BWP7T $T=180160 412000 1 180 $X=178190 $Y=411765
X1132 309 1 2 928 INVD1BWP7T $T=181280 404160 0 0 $X=180990 $Y=403925
X1133 964 1 2 277 INVD1BWP7T $T=184640 396320 0 180 $X=182670 $Y=392110
X1134 316 1 2 949 INVD1BWP7T $T=185760 412000 0 0 $X=185470 $Y=411765
X1135 931 1 2 981 INVD1BWP7T $T=186320 388480 1 0 $X=186030 $Y=384270
X1136 329 1 2 948 INVD1BWP7T $T=190800 380640 0 180 $X=188830 $Y=376430
X1137 334 1 2 994 INVD1BWP7T $T=195280 364960 1 180 $X=193310 $Y=364725
X1138 971 1 2 346 INVD1BWP7T $T=208160 412000 0 180 $X=206190 $Y=407790
X1139 972 1 2 1009 INVD1BWP7T $T=209280 388480 1 0 $X=208990 $Y=384270
X1140 1002 1 2 1001 INVD1BWP7T $T=213200 372800 0 180 $X=211230 $Y=368590
X1141 984 1 2 356 INVD1BWP7T $T=212080 380640 0 0 $X=211790 $Y=380405
X1142 965 1 2 1004 INVD1BWP7T $T=213200 388480 0 0 $X=212910 $Y=388245
X1143 1016 1 2 992 INVD1BWP7T $T=221600 380640 1 180 $X=219630 $Y=380405
X1144 385 1 2 381 INVD1BWP7T $T=237840 404160 1 180 $X=235870 $Y=403925
X1145 448 1 2 447 INVD1BWP7T $T=292720 380640 0 180 $X=290750 $Y=376430
X1146 451 1 2 450 INVD1BWP7T $T=295520 357120 1 180 $X=293550 $Y=356885
X1147 465 1 2 460 INVD1BWP7T $T=300560 380640 0 180 $X=298590 $Y=376430
X1148 530 1 2 1063 INVD1BWP7T $T=353760 412000 0 180 $X=351790 $Y=407790
X1149 592 1 2 584 INVD1BWP7T $T=406400 412000 0 180 $X=404430 $Y=407790
X1150 1 2 ICV_14 $T=59760 396320 1 0 $X=59470 $Y=392110
X1151 1 2 ICV_14 $T=138720 396320 0 0 $X=138430 $Y=396085
X1152 1 2 ICV_14 $T=196400 380640 0 0 $X=196110 $Y=380405
X1153 1 2 ICV_14 $T=213200 372800 1 0 $X=212910 $Y=368590
X1154 1 2 ICV_14 $T=238400 364960 0 0 $X=238110 $Y=364725
X1155 1 2 ICV_14 $T=254080 412000 0 0 $X=253790 $Y=411765
X1156 1 2 ICV_14 $T=263040 412000 1 0 $X=262750 $Y=407790
X1157 1 2 ICV_14 $T=270880 388480 0 0 $X=270590 $Y=388245
X1158 1 2 ICV_14 $T=280400 372800 1 0 $X=280110 $Y=368590
X1159 1 2 ICV_14 $T=280400 372800 0 0 $X=280110 $Y=372565
X1160 1 2 ICV_14 $T=349280 380640 0 0 $X=348990 $Y=380405
X1161 1 2 ICV_14 $T=364400 404160 1 0 $X=364110 $Y=399950
X1162 1 2 ICV_14 $T=371120 357120 0 0 $X=370830 $Y=356885
X1163 1 2 ICV_14 $T=392400 364960 1 0 $X=392110 $Y=360750
X1164 1 2 ICV_14 $T=399120 412000 1 0 $X=398830 $Y=407790
X1165 1 2 ICV_14 $T=401360 396320 0 0 $X=401070 $Y=396085
X1166 1 2 ICV_14 $T=406400 404160 0 0 $X=406110 $Y=403925
X1167 1 2 ICV_14 $T=448400 404160 0 0 $X=448110 $Y=403925
X1168 1 2 ICV_14 $T=448400 412000 1 0 $X=448110 $Y=407790
X1169 1026 389 1 2 BUFFD2BWP7T $T=233920 380640 1 180 $X=230270 $Y=380405
X1170 1030 373 1 2 BUFFD2BWP7T $T=238400 364960 1 180 $X=234750 $Y=364725
X1171 1173 565 1 2 BUFFD2BWP7T $T=460160 364960 0 0 $X=459870 $Y=364725
X1172 648 474 1 2 BUFFD2BWP7T $T=463520 388480 1 180 $X=459870 $Y=388245
X1173 436 631 532 617 1 2 DFCNQD2BWP7T $T=448400 412000 0 180 $X=435230 $Y=407790
X1174 1 2 DCAP16BWP7T $T=128080 412000 0 0 $X=127790 $Y=411765
X1175 1 2 DCAP16BWP7T $T=231680 388480 0 0 $X=231390 $Y=388245
X1176 1 2 DCAP16BWP7T $T=235040 357120 0 0 $X=234750 $Y=356885
X1177 1 2 DCAP16BWP7T $T=245120 372800 0 0 $X=244830 $Y=372565
X1178 1 2 DCAP16BWP7T $T=245120 412000 0 0 $X=244830 $Y=411765
X1179 1 2 DCAP16BWP7T $T=261360 388480 1 0 $X=261070 $Y=384270
X1180 1 2 DCAP16BWP7T $T=287120 364960 1 0 $X=286830 $Y=360750
X1181 1 2 DCAP16BWP7T $T=287120 388480 1 0 $X=286830 $Y=384270
X1182 1 2 DCAP16BWP7T $T=298320 372800 1 0 $X=298030 $Y=368590
X1183 1 2 DCAP16BWP7T $T=305040 388480 0 0 $X=304750 $Y=388245
X1184 1 2 DCAP16BWP7T $T=307840 364960 0 0 $X=307550 $Y=364725
X1185 1 2 DCAP16BWP7T $T=316240 364960 1 0 $X=315950 $Y=360750
X1186 1 2 DCAP16BWP7T $T=329120 412000 0 0 $X=328830 $Y=411765
X1187 1 2 DCAP16BWP7T $T=339760 404160 0 0 $X=339470 $Y=403925
X1188 1 2 DCAP16BWP7T $T=343680 364960 1 0 $X=343390 $Y=360750
X1189 1 2 DCAP16BWP7T $T=352640 404160 0 0 $X=352350 $Y=403925
X1190 1 2 DCAP16BWP7T $T=358800 388480 1 0 $X=358510 $Y=384270
X1191 1 2 DCAP16BWP7T $T=360480 357120 0 0 $X=360190 $Y=356885
X1192 1 2 DCAP16BWP7T $T=371120 380640 0 0 $X=370830 $Y=380405
X1193 1 2 DCAP16BWP7T $T=371120 404160 0 0 $X=370830 $Y=403925
X1194 1 2 DCAP16BWP7T $T=376160 372800 0 0 $X=375870 $Y=372565
X1195 1 2 DCAP16BWP7T $T=383440 412000 0 0 $X=383150 $Y=411765
X1196 1 2 DCAP16BWP7T $T=385120 388480 0 0 $X=384830 $Y=388245
X1197 1 2 DCAP16BWP7T $T=386800 380640 0 0 $X=386510 $Y=380405
X1198 1 2 DCAP16BWP7T $T=387360 404160 1 0 $X=387070 $Y=399950
X1199 1 2 DCAP16BWP7T $T=390720 364960 0 0 $X=390430 $Y=364725
X1200 1 2 DCAP16BWP7T $T=401360 404160 1 0 $X=401070 $Y=399950
X1201 1 2 DCAP16BWP7T $T=413120 364960 1 0 $X=412830 $Y=360750
X1202 1 2 DCAP16BWP7T $T=413120 396320 0 0 $X=412830 $Y=396085
X1203 1 2 DCAP16BWP7T $T=413120 404160 0 0 $X=412830 $Y=403925
X1204 1 2 DCAP16BWP7T $T=425440 404160 0 0 $X=425150 $Y=403925
X1205 1 2 DCAP16BWP7T $T=427680 404160 1 0 $X=427390 $Y=399950
X1206 1 2 DCAP16BWP7T $T=432720 388480 0 0 $X=432430 $Y=388245
X1207 1 2 DCAP16BWP7T $T=435520 412000 0 0 $X=435230 $Y=411765
X1208 1 2 DCAP16BWP7T $T=436080 380640 1 0 $X=435790 $Y=376430
X1209 1 2 DCAP16BWP7T $T=441120 396320 0 0 $X=440830 $Y=396085
X1210 1 2 DCAP16BWP7T $T=455120 380640 1 0 $X=454830 $Y=376430
X1211 1 2 DCAP16BWP7T $T=455120 396320 0 0 $X=454830 $Y=396085
X1212 796 1 2 17 CKND1BWP7T $T=24480 380640 0 0 $X=24190 $Y=380405
X1213 795 1 2 112 CKND1BWP7T $T=67040 396320 0 180 $X=65070 $Y=392110
X1214 55 1 2 109 CKND1BWP7T $T=71520 412000 1 180 $X=69550 $Y=411765
X1215 95 1 2 133 CKND1BWP7T $T=71520 404160 0 0 $X=71230 $Y=403925
X1216 97 1 2 857 CKND1BWP7T $T=88880 388480 1 180 $X=86910 $Y=388245
X1217 811 1 2 189 CKND1BWP7T $T=102320 412000 1 0 $X=102030 $Y=407790
X1218 142 1 2 920 CKND1BWP7T $T=146000 364960 0 180 $X=144030 $Y=360750
X1219 245 1 2 940 CKND1BWP7T $T=166160 388480 0 180 $X=164190 $Y=384270
X1220 956 1 2 959 CKND1BWP7T $T=178480 380640 0 180 $X=176510 $Y=376430
X1221 998 1 2 1007 CKND1BWP7T $T=221040 396320 1 180 $X=219070 $Y=396085
X1222 440 1 2 437 CKND1BWP7T $T=279840 364960 0 180 $X=277870 $Y=360750
X1223 527 1 2 1072 CKND1BWP7T $T=351520 412000 0 180 $X=349550 $Y=407790
X1224 1122 586 1 2 INVD4BWP7T $T=397440 404160 1 0 $X=397150 $Y=399950
X1225 368 1 2 355 BUFFD3BWP7T $T=216560 357120 1 180 $X=212350 $Y=356885
X1226 1029 1 2 393 BUFFD3BWP7T $T=236720 372800 1 180 $X=232510 $Y=372565
X1227 430 1 2 411 BUFFD3BWP7T $T=272560 412000 0 180 $X=268350 $Y=407790
X1228 421 1 2 522 BUFFD3BWP7T $T=337520 412000 1 0 $X=337230 $Y=407790
X1229 1169 1168 609 1 2 CKXOR2D4BWP7T $T=441120 396320 1 180 $X=428510 $Y=396085
X1230 385 398 2 381 1 395 1021 AOI22D1BWP7T $T=237840 412000 1 180 $X=233630 $Y=411765
X1231 1056 446 2 1059 1 1046 1067 AOI22D1BWP7T $T=294960 372800 1 180 $X=290750 $Y=372565
X1232 466 498 2 464 1 469 497 AOI22D1BWP7T $T=317920 372800 1 0 $X=317630 $Y=368590
X1233 1060 534 2 1109 1 528 1113 AOI22D1BWP7T $T=354880 380640 0 0 $X=354590 $Y=380405
X1234 466 538 2 464 1 551 1128 AOI22D1BWP7T $T=373920 364960 0 0 $X=373630 $Y=364725
X1235 563 561 2 557 1 1129 554 AOI22D1BWP7T $T=381760 388480 0 180 $X=377550 $Y=384270
X1236 594 591 2 1152 1 579 1141 AOI22D1BWP7T $T=407520 372800 1 180 $X=403310 $Y=372565
X1237 1161 591 2 599 1 579 1159 AOI22D1BWP7T $T=422640 380640 1 180 $X=418430 $Y=380405
X1238 563 606 2 557 1 1150 598 AOI22D1BWP7T $T=442800 357120 1 180 $X=438590 $Y=356885
X1239 563 597 2 557 1 1170 627 AOI22D1BWP7T $T=443360 380640 0 0 $X=443070 $Y=380405
X1240 563 1168 2 557 1 633 624 AOI22D1BWP7T $T=443920 388480 0 0 $X=443630 $Y=388245
X1241 933 1017 2 1019 371 1 OAI21D1BWP7T $T=220480 412000 1 0 $X=220190 $Y=407790
X1242 409 1038 2 425 1045 1 OAI21D1BWP7T $T=266400 380640 1 0 $X=266110 $Y=376430
X1243 493 1075 2 489 492 1 OAI21D1BWP7T $T=317360 404160 0 180 $X=313710 $Y=399950
X1244 493 1084 2 501 496 1 OAI21D1BWP7T $T=317360 404160 0 0 $X=317070 $Y=403925
X1245 556 1166 2 1156 1169 1 OAI21D1BWP7T $T=433840 380640 1 180 $X=430190 $Y=380405
X1246 401 2 391 1 CKND12BWP7T $T=237840 364960 0 180 $X=228590 $Y=360750
X1247 857 2 19 859 1 NR2D4BWP7T $T=104560 396320 0 0 $X=104270 $Y=396085
X1248 235 2 245 243 1 NR2D4BWP7T $T=146000 380640 0 0 $X=145710 $Y=380405
X1249 77 823 2 1 INVD2BWP7T $T=53600 404160 0 180 $X=51070 $Y=399950
X1250 130 797 2 1 INVD2BWP7T $T=73200 372800 1 180 $X=70670 $Y=372565
X1251 137 126 2 1 INVD2BWP7T $T=73200 380640 0 180 $X=70670 $Y=376430
X1252 850 173 2 1 INVD2BWP7T $T=92240 396320 1 0 $X=91950 $Y=392110
X1253 872 76 2 1 INVD2BWP7T $T=98400 372800 0 0 $X=98110 $Y=372565
X1254 908 831 2 1 INVD2BWP7T $T=128640 388480 1 180 $X=126110 $Y=388245
X1255 211 806 2 1 INVD2BWP7T $T=133120 388480 0 180 $X=130590 $Y=384270
X1256 818 897 2 1 INVD2BWP7T $T=133680 396320 1 0 $X=133390 $Y=392110
X1257 910 73 2 1 INVD2BWP7T $T=144320 388480 0 180 $X=141790 $Y=384270
X1258 939 235 2 1 INVD2BWP7T $T=154960 380640 1 180 $X=152430 $Y=380405
X1259 932 933 2 1 INVD2BWP7T $T=157200 396320 0 180 $X=154670 $Y=392110
X1260 953 990 2 1 INVD2BWP7T $T=190240 364960 0 0 $X=189950 $Y=364725
X1261 999 993 2 1 INVD2BWP7T $T=205920 364960 0 0 $X=205630 $Y=364725
X1262 445 444 2 1 INVD2BWP7T $T=289920 357120 0 0 $X=289630 $Y=356885
X1263 379 512 2 1 INVD2BWP7T $T=334720 372800 0 0 $X=334430 $Y=372565
X1264 495 505 2 1 INVD2BWP7T $T=347040 380640 0 0 $X=346750 $Y=380405
X1265 526 525 2 1 INVD2BWP7T $T=352080 388480 1 180 $X=349550 $Y=388245
X1266 538 523 2 1 INVD2BWP7T $T=384000 372800 1 0 $X=383710 $Y=368590
X1267 570 511 2 1 INVD2BWP7T $T=399120 396320 0 0 $X=398830 $Y=396085
X1268 1168 610 2 1 INVD2BWP7T $T=432720 388480 1 180 $X=430190 $Y=388245
X1269 1052 528 1 2 1107 CKXOR2D1BWP7T $T=348160 380640 1 0 $X=347870 $Y=376430
X1270 581 579 1 2 1148 CKXOR2D1BWP7T $T=396880 357120 0 0 $X=396590 $Y=356885
X1271 1148 1150 1 2 1144 CKXOR2D1BWP7T $T=400800 364960 0 0 $X=400510 $Y=364725
X1272 389 383 871 1 2 CKXOR2D2BWP7T $T=232800 364960 1 180 $X=226350 $Y=364725
X1273 411 403 883 1 2 CKXOR2D2BWP7T $T=255760 388480 1 180 $X=249310 $Y=388245
X1274 566 1130 552 1 2 CKXOR2D2BWP7T $T=383440 412000 1 180 $X=376990 $Y=411765
X1275 570 1131 562 1 2 CKXOR2D2BWP7T $T=386800 380640 1 180 $X=380350 $Y=380405
X1276 589 585 334 1 2 CKXOR2D2BWP7T $T=403040 412000 1 180 $X=396590 $Y=411765
X1277 2 1 DCAP32BWP7T $T=130880 404160 0 0 $X=130590 $Y=403925
X1278 2 1 DCAP32BWP7T $T=225520 372800 1 0 $X=225230 $Y=368590
X1279 396 1 2 380 BUFFD5BWP7T $T=235600 380640 0 180 $X=229150 $Y=376430
X1280 520 1 2 404 BUFFD5BWP7T $T=340320 412000 0 0 $X=340030 $Y=411765
X1281 1073 1087 500 503 1 2 OAI21D0BWP7T $T=319040 404160 1 0 $X=318750 $Y=399950
X1282 1049 1088 1081 509 1 2 OAI21D0BWP7T $T=321840 372800 0 0 $X=321550 $Y=372565
X1283 1093 1095 515 503 1 2 OAI21D0BWP7T $T=334160 404160 0 0 $X=333870 $Y=403925
X1284 1098 1105 529 509 1 2 OAI21D0BWP7T $T=350960 396320 0 0 $X=350670 $Y=396085
X1285 1114 1117 539 509 1 2 OAI21D0BWP7T $T=361600 404160 1 0 $X=361310 $Y=399950
X1286 1116 1123 550 1125 1 2 OAI21D0BWP7T $T=374480 380640 1 0 $X=374190 $Y=376430
X1287 1133 1131 556 1126 1 2 OAI21D0BWP7T $T=380640 372800 0 180 $X=377550 $Y=368590
X1288 583 1151 580 1140 1 2 OAI21D0BWP7T $T=405840 388480 0 180 $X=402750 $Y=384270
X1289 1145 1158 596 509 1 2 OAI21D0BWP7T $T=420400 364960 1 180 $X=417310 $Y=364725
X1290 1154 1160 601 509 1 2 OAI21D0BWP7T $T=423200 396320 0 180 $X=420110 $Y=392110
X1291 1159 1146 602 1162 1 2 OAI21D0BWP7T $T=421520 388480 1 0 $X=421230 $Y=384270
X1292 399 1025 1022 1021 376 1 2 XNR4D0BWP7T $T=237840 396320 1 180 $X=224670 $Y=396085
X1293 1023 1024 386 382 375 1 2 XNR4D2BWP7T $T=237840 404160 0 180 $X=224110 $Y=399950
X1294 1023 1028 388 387 378 1 2 XNR4D2BWP7T $T=238960 412000 0 180 $X=225230 $Y=407790
X1295 419 1036 410 1021 387 1 2 XNR4D2BWP7T $T=263040 412000 0 180 $X=249310 $Y=407790
X1296 428 1047 421 420 417 1 2 XNR4D2BWP7T $T=273120 412000 1 180 $X=259390 $Y=411765
X1297 381 942 385 1 2 390 MUX2ND1BWP7T $T=225520 388480 0 0 $X=225230 $Y=388245
X1298 381 950 385 1 2 397 MUX2ND1BWP7T $T=229440 396320 1 0 $X=229150 $Y=392110
X1299 519 521 517 1 2 513 MUX2ND1BWP7T $T=342000 357120 1 180 $X=335550 $Y=356885
X1300 369 363 1 2 1014 XNR2D1BWP7T $T=221600 364960 1 180 $X=216270 $Y=364725
X1301 379 1020 1 2 1018 XNR2D1BWP7T $T=227760 380640 1 180 $X=222430 $Y=380405
X1302 379 1020 1 2 983 XNR2D1BWP7T $T=228880 372800 1 180 $X=223550 $Y=372565
X1303 577 505 1 2 1112 XNR2D1BWP7T $T=393520 380640 0 180 $X=388190 $Y=376430
X1304 579 1100 1 2 1138 XNR2D1BWP7T $T=397440 372800 1 180 $X=392110 $Y=372565
X1305 78 15 2 1 CKND2BWP7T $T=53600 404160 1 180 $X=51070 $Y=403925
X1306 944 1 2 930 CKND0BWP7T $T=165600 380640 0 180 $X=163630 $Y=376430
X1307 256 1 2 961 CKND0BWP7T $T=184080 380640 0 0 $X=183790 $Y=380405
X1308 333 1 2 915 CKND0BWP7T $T=191920 404160 1 0 $X=191630 $Y=399950
X1309 469 1 2 453 CKND0BWP7T $T=304480 357120 1 180 $X=302510 $Y=356885
X1310 524 1 2 1065 CKND0BWP7T $T=347040 412000 0 180 $X=345070 $Y=407790
X1311 377 384 1 2 1023 CKXOR2D0BWP7T $T=224960 412000 0 0 $X=224670 $Y=411765
X1312 1044 2 422 1049 1046 424 1 AOI22D2BWP7T $T=264160 372800 1 0 $X=263870 $Y=368590
X1313 1086 2 505 1079 495 1083 1 AOI22D2BWP7T $T=322960 388480 1 180 $X=315950 $Y=388245
X1314 466 2 445 507 440 464 1 AOI22D2BWP7T $T=316800 364960 0 0 $X=316510 $Y=364725
X1315 1092 2 505 1098 495 1094 1 AOI22D2BWP7T $T=338080 388480 0 0 $X=337790 $Y=388245
X1316 1111 2 534 1116 528 1099 1 AOI22D2BWP7T $T=356000 372800 0 0 $X=355710 $Y=372565
X1317 563 2 565 572 569 557 1 AOI22D2BWP7T $T=381760 357120 0 0 $X=381470 $Y=356885
X1318 1027 385 381 1024 1 2 MUX2ND0BWP7T $T=236160 404160 1 180 $X=231390 $Y=403925
X1319 1107 571 1136 1133 1 2 MUX2ND0BWP7T $T=386240 364960 0 0 $X=385950 $Y=364725
X1320 1112 578 584 1137 1 2 MUX2ND0BWP7T $T=394640 412000 1 0 $X=394350 $Y=407790
X1321 1138 633 622 1166 1 2 MUX2ND0BWP7T $T=449520 372800 1 180 $X=444750 $Y=372565
X1322 379 1074 471 466 464 2 1 AOI22D0BWP7T $T=307840 364960 1 180 $X=304190 $Y=364725
X1323 119 1 2 156 CKBD0BWP7T $T=84400 357120 0 0 $X=84110 $Y=356885
X1324 939 951 274 923 2 1 271 AO211D1BWP7T $T=170640 380640 1 180 $X=165870 $Y=380405
X1325 122 2 845 816 1 NR2D1BWP7T $T=69280 396320 0 180 $X=66750 $Y=392110
X1326 149 2 850 859 1 NR2D1BWP7T $T=84400 396320 1 0 $X=84110 $Y=392110
X1327 823 2 158 150 1 NR2D1BWP7T $T=91680 404160 0 180 $X=89150 $Y=399950
X1328 130 2 163 872 1 NR2D1BWP7T $T=93920 372800 1 0 $X=93630 $Y=368590
X1329 823 2 179 55 1 NR2D1BWP7T $T=95600 412000 0 0 $X=95310 $Y=411765
X1330 872 2 882 19 1 NR2D1BWP7T $T=104560 388480 1 0 $X=104270 $Y=384270
X1331 887 2 901 906 1 NR2D1BWP7T $T=123600 412000 1 0 $X=123310 $Y=407790
X1332 914 2 894 227 1 NR2D1BWP7T $T=144320 364960 0 180 $X=141790 $Y=360750
X1333 232 2 921 925 1 NR2D1BWP7T $T=144320 404160 1 0 $X=144030 $Y=399950
X1334 237 2 247 931 1 NR2D1BWP7T $T=150480 396320 1 0 $X=150190 $Y=392110
X1335 929 2 923 256 1 NR2D1BWP7T $T=168400 388480 0 180 $X=165870 $Y=384270
X1336 297 2 957 287 1 NR2D1BWP7T $T=174560 412000 1 180 $X=172030 $Y=411765
X1337 967 2 254 273 1 NR2D1BWP7T $T=178480 404160 1 180 $X=175950 $Y=403925
X1338 305 2 307 287 1 NR2D1BWP7T $T=183520 412000 0 180 $X=180990 $Y=407790
X1339 317 2 309 977 1 NR2D1BWP7T $T=185760 404160 1 180 $X=183230 $Y=403925
X1340 329 2 977 933 1 NR2D1BWP7T $T=194160 396320 1 180 $X=191630 $Y=396085
X1341 934 2 996 1002 1 NR2D1BWP7T $T=199200 396320 1 180 $X=196670 $Y=396085
X1342 329 2 344 239 1 NR2D1BWP7T $T=196960 412000 0 0 $X=196670 $Y=411765
X1343 263 2 347 1006 1 NR2D1BWP7T $T=205920 372800 0 0 $X=205630 $Y=372565
X1344 958 2 349 988 1 NR2D1BWP7T $T=207040 404160 1 0 $X=206750 $Y=399950
X1345 1014 2 1016 334 1 NR2D1BWP7T $T=219360 380640 0 180 $X=216830 $Y=376430
X1346 1073 1080 500 1087 1 2 AOI21D0BWP7T $T=318480 396320 0 0 $X=318190 $Y=396085
X1347 1049 1078 1081 1088 1 2 AOI21D0BWP7T $T=320160 380640 1 0 $X=319870 $Y=376430
X1348 1093 1096 515 1095 1 2 AOI21D0BWP7T $T=336960 404160 0 0 $X=336670 $Y=403925
X1349 1114 1115 539 1117 1 2 AOI21D0BWP7T $T=358800 396320 1 0 $X=358510 $Y=392110
X1350 1116 1125 550 556 1 2 AOI21D0BWP7T $T=380640 380640 1 0 $X=380350 $Y=376430
X1351 583 1140 580 556 1 2 AOI21D0BWP7T $T=398560 388480 0 180 $X=395470 $Y=384270
X1352 1154 1163 601 1160 1 2 AOI21D0BWP7T $T=428240 396320 1 0 $X=427950 $Y=392110
X1353 1159 1162 612 556 1 2 AOI21D0BWP7T $T=431040 388480 1 0 $X=430750 $Y=384270
X1354 32 794 21 793 2 1 798 NR4D1BWP7T $T=30640 364960 1 180 $X=24750 $Y=364725
X1355 54 810 792 23 2 1 807 NR4D1BWP7T $T=44080 364960 1 180 $X=38190 $Y=364725
X1356 51 814 816 820 2 1 819 NR4D1BWP7T $T=43520 396320 0 0 $X=43230 $Y=396085
X1357 75 827 817 83 2 1 84 NR4D1BWP7T $T=50800 412000 0 0 $X=50510 $Y=411765
X1358 110 840 839 101 2 1 98 NR4D1BWP7T $T=65920 357120 1 180 $X=60030 $Y=356885
X1359 146 816 820 49 2 1 136 NR4D1BWP7T $T=85520 364960 0 180 $X=79630 $Y=360750
X1360 855 856 802 844 2 1 11 NR4D1BWP7T $T=83280 380640 1 0 $X=82990 $Y=376430
X1361 170 841 866 870 2 1 173 NR4D1BWP7T $T=91680 388480 0 0 $X=91390 $Y=388245
X1362 175 811 158 172 2 1 116 NR4D1BWP7T $T=97840 404160 1 180 $X=91950 $Y=403925
X1363 873 63 101 867 2 1 869 NR4D1BWP7T $T=100080 364960 1 180 $X=94190 $Y=364725
X1364 209 814 56 853 2 1 889 NR4D1BWP7T $T=115200 372800 0 180 $X=109310 $Y=368590
X1365 218 841 214 876 2 1 902 NR4D1BWP7T $T=128640 388480 0 180 $X=122750 $Y=384270
X1366 937 260 255 243 2 1 237 NR4D1BWP7T $T=156640 388480 0 180 $X=150750 $Y=384270
X1367 955 277 276 271 2 1 267 NR4D1BWP7T $T=170640 404160 1 180 $X=164750 $Y=403925
X1368 936 260 949 282 2 1 938 NR4D1BWP7T $T=165600 412000 1 0 $X=165310 $Y=407790
X1369 924 299 949 304 2 1 287 NR4D1BWP7T $T=175680 412000 1 0 $X=175390 $Y=407790
X1370 352 260 346 353 2 1 305 NR4D1BWP7T $T=206480 412000 0 0 $X=206190 $Y=411765
X1371 351 287 305 1013 2 1 323 NR4D1BWP7T $T=209840 412000 1 0 $X=209550 $Y=407790
X1372 804 803 25 801 2 1 796 OR4D1BWP7T $T=30640 380640 1 180 $X=25870 $Y=380405
X1373 277 2 284 940 961 1 AOI21D2BWP7T $T=170080 396320 1 0 $X=169790 $Y=392110
X1374 239 2 317 329 263 1 AOI21D2BWP7T $T=194160 404160 0 0 $X=193870 $Y=403925
X1375 8 1 791 9 2 ND2D1BWP7T $T=22800 372800 1 0 $X=22510 $Y=368590
X1376 27 1 31 806 2 ND2D1BWP7T $T=28960 357120 0 0 $X=28670 $Y=356885
X1377 27 1 37 809 2 ND2D1BWP7T $T=37920 372800 0 0 $X=37630 $Y=372565
X1378 37 1 808 22 2 ND2D1BWP7T $T=40160 388480 1 180 $X=37630 $Y=388245
X1379 43 1 807 39 2 ND2D1BWP7T $T=41280 357120 0 0 $X=40990 $Y=356885
X1380 14 1 39 818 2 ND2D1BWP7T $T=42960 364960 1 0 $X=42670 $Y=360750
X1381 8 1 44 14 2 ND2D1BWP7T $T=43520 357120 0 0 $X=43230 $Y=356885
X1382 815 1 60 52 2 ND2D1BWP7T $T=48000 412000 1 180 $X=45470 $Y=411765
X1383 5 1 790 73 2 ND2D1BWP7T $T=53600 372800 1 180 $X=51070 $Y=372565
X1384 806 1 79 818 2 ND2D1BWP7T $T=51920 364960 1 0 $X=51630 $Y=360750
X1385 8 1 43 831 2 ND2D1BWP7T $T=52480 357120 0 0 $X=52190 $Y=356885
X1386 809 1 74 76 2 ND2D1BWP7T $T=55280 364960 1 180 $X=52750 $Y=364725
X1387 5 1 68 809 2 ND2D1BWP7T $T=53600 372800 0 0 $X=53310 $Y=372565
X1388 8 1 80 809 2 ND2D1BWP7T $T=54160 364960 1 0 $X=53870 $Y=360750
X1389 68 1 829 833 2 ND2D1BWP7T $T=54720 380640 1 0 $X=54430 $Y=376430
X1390 831 1 69 76 2 ND2D1BWP7T $T=55280 372800 1 0 $X=54990 $Y=368590
X1391 818 1 825 809 2 ND2D1BWP7T $T=58080 364960 1 180 $X=55550 $Y=364725
X1392 831 1 833 5 2 ND2D1BWP7T $T=59200 372800 1 180 $X=56670 $Y=372565
X1393 806 1 72 97 2 ND2D1BWP7T $T=58080 364960 0 0 $X=57790 $Y=364725
X1394 73 1 788 97 2 ND2D1BWP7T $T=58640 380640 1 0 $X=58350 $Y=376430
X1395 806 1 94 91 2 ND2D1BWP7T $T=61440 372800 1 180 $X=58910 $Y=372565
X1396 77 1 88 96 2 ND2D1BWP7T $T=62000 412000 1 180 $X=59470 $Y=411765
X1397 36 1 102 788 2 ND2D1BWP7T $T=62560 364960 0 180 $X=60030 $Y=360750
X1398 790 1 838 28 2 ND2D1BWP7T $T=61440 372800 0 0 $X=61150 $Y=372565
X1399 109 1 106 815 2 ND2D1BWP7T $T=64240 412000 1 180 $X=61710 $Y=411765
X1400 72 1 842 825 2 ND2D1BWP7T $T=63120 364960 0 0 $X=62830 $Y=364725
X1401 117 1 839 36 2 ND2D1BWP7T $T=65920 364960 0 180 $X=63390 $Y=360750
X1402 806 1 104 76 2 ND2D1BWP7T $T=63680 372800 0 0 $X=63390 $Y=372565
X1403 79 1 844 81 2 ND2D1BWP7T $T=64240 372800 1 0 $X=63950 $Y=368590
X1404 57 1 840 845 2 ND2D1BWP7T $T=65920 372800 0 0 $X=65630 $Y=372565
X1405 46 1 123 109 2 ND2D1BWP7T $T=67600 412000 0 0 $X=67310 $Y=411765
X1406 121 1 847 112 2 ND2D1BWP7T $T=70400 388480 1 180 $X=67870 $Y=388245
X1407 797 1 121 848 2 ND2D1BWP7T $T=68720 372800 0 0 $X=68430 $Y=372565
X1408 837 1 125 114 2 ND2D1BWP7T $T=69280 404160 0 0 $X=68990 $Y=403925
X1409 22 1 851 44 2 ND2D1BWP7T $T=70960 388480 0 0 $X=70670 $Y=388245
X1410 849 1 137 831 2 ND2D1BWP7T $T=79920 380640 0 0 $X=79630 $Y=380405
X1411 831 1 160 97 2 ND2D1BWP7T $T=87200 388480 1 0 $X=86910 $Y=384270
X1412 806 1 862 5 2 ND2D1BWP7T $T=91120 380640 0 180 $X=88590 $Y=376430
X1413 868 1 98 862 2 ND2D1BWP7T $T=93360 380640 0 180 $X=90830 $Y=376430
X1414 68 1 867 862 2 ND2D1BWP7T $T=93920 364960 1 180 $X=91390 $Y=364725
X1415 78 1 176 815 2 ND2D1BWP7T $T=92240 412000 0 0 $X=91950 $Y=411765
X1416 76 1 865 73 2 ND2D1BWP7T $T=96160 372800 0 0 $X=95870 $Y=372565
X1417 143 1 180 877 2 ND2D1BWP7T $T=97840 412000 0 0 $X=97550 $Y=411765
X1418 187 1 182 76 2 ND2D1BWP7T $T=102880 357120 1 180 $X=100350 $Y=356885
X1419 824 1 192 888 2 ND2D1BWP7T $T=101760 380640 0 0 $X=101470 $Y=380405
X1420 849 1 169 806 2 ND2D1BWP7T $T=108480 380640 0 180 $X=105950 $Y=376430
X1421 27 1 868 831 2 ND2D1BWP7T $T=111840 388480 0 180 $X=109310 $Y=384270
X1422 806 1 893 843 2 ND2D1BWP7T $T=112400 380640 1 180 $X=109870 $Y=380405
X1423 906 1 202 907 2 ND2D1BWP7T $T=128640 412000 0 180 $X=126110 $Y=407790
X1424 117 1 909 104 2 ND2D1BWP7T $T=129760 357120 0 0 $X=129470 $Y=356885
X1425 906 1 861 883 2 ND2D1BWP7T $T=134240 404160 0 180 $X=131710 $Y=399950
X1426 14 1 167 5 2 ND2D1BWP7T $T=134240 372800 0 0 $X=133950 $Y=372565
X1427 849 1 895 14 2 ND2D1BWP7T $T=135920 357120 0 0 $X=135630 $Y=356885
X1428 27 1 904 73 2 ND2D1BWP7T $T=140400 388480 0 180 $X=137870 $Y=384270
X1429 843 1 872 226 2 ND2D1BWP7T $T=140960 380640 0 180 $X=138430 $Y=376430
X1430 142 1 900 914 2 ND2D1BWP7T $T=139840 364960 1 0 $X=139550 $Y=360750
X1431 230 1 908 225 2 ND2D1BWP7T $T=143760 357120 1 180 $X=141230 $Y=356885
X1432 236 1 918 920 2 ND2D1BWP7T $T=148800 372800 1 180 $X=146270 $Y=372565
X1433 246 1 881 241 2 ND2D1BWP7T $T=152160 357120 1 180 $X=149630 $Y=356885
X1434 241 1 863 234 2 ND2D1BWP7T $T=153840 364960 0 180 $X=151310 $Y=360750
X1435 935 1 240 932 2 ND2D1BWP7T $T=154960 396320 0 180 $X=152430 $Y=392110
X1436 939 1 268 944 2 ND2D1BWP7T $T=163920 380640 0 0 $X=163630 $Y=380405
X1437 940 1 262 947 2 ND2D1BWP7T $T=164480 388480 0 0 $X=164190 $Y=388245
X1438 935 1 945 940 2 ND2D1BWP7T $T=164480 396320 0 0 $X=164190 $Y=396085
X1439 940 1 258 948 2 ND2D1BWP7T $T=165040 396320 1 0 $X=164750 $Y=392110
X1440 944 1 275 947 2 ND2D1BWP7T $T=166720 388480 0 0 $X=166430 $Y=388245
X1441 944 1 278 953 2 ND2D1BWP7T $T=167840 372800 1 0 $X=167550 $Y=368590
X1442 944 1 280 948 2 ND2D1BWP7T $T=168960 388480 0 0 $X=168670 $Y=388245
X1443 954 1 289 947 2 ND2D1BWP7T $T=170640 380640 0 0 $X=170350 $Y=380405
X1444 957 1 253 916 2 ND2D1BWP7T $T=173440 412000 0 180 $X=170910 $Y=407790
X1445 959 1 922 947 2 ND2D1BWP7T $T=174000 372800 0 180 $X=171470 $Y=368590
X1446 954 1 290 935 2 ND2D1BWP7T $T=175120 396320 1 180 $X=172590 $Y=396085
X1447 939 1 296 959 2 ND2D1BWP7T $T=174000 364960 1 0 $X=173710 $Y=360750
X1448 959 1 286 953 2 ND2D1BWP7T $T=176240 372800 0 180 $X=173710 $Y=368590
X1449 959 1 288 948 2 ND2D1BWP7T $T=176800 380640 0 180 $X=174270 $Y=376430
X1450 289 1 927 966 2 ND2D1BWP7T $T=175120 380640 0 0 $X=174830 $Y=380405
X1451 935 1 964 944 2 ND2D1BWP7T $T=175120 388480 0 0 $X=174830 $Y=388245
X1452 963 1 294 935 2 ND2D1BWP7T $T=177360 396320 1 180 $X=174830 $Y=396085
X1453 965 1 269 944 2 ND2D1BWP7T $T=177920 404160 0 180 $X=175390 $Y=399950
X1454 954 1 303 948 2 ND2D1BWP7T $T=177360 388480 0 0 $X=177070 $Y=388245
X1455 963 1 261 965 2 ND2D1BWP7T $T=177360 396320 0 0 $X=177070 $Y=396085
X1456 973 1 969 959 2 ND2D1BWP7T $T=180160 372800 1 180 $X=177630 $Y=372565
X1457 939 1 283 972 2 ND2D1BWP7T $T=178480 364960 1 0 $X=178190 $Y=360750
X1458 973 1 293 963 2 ND2D1BWP7T $T=180720 396320 0 180 $X=178190 $Y=392110
X1459 954 1 311 965 2 ND2D1BWP7T $T=179600 396320 0 0 $X=179310 $Y=396085
X1460 973 1 300 932 2 ND2D1BWP7T $T=180160 388480 0 0 $X=179870 $Y=388245
X1461 972 1 308 953 2 ND2D1BWP7T $T=182960 364960 0 180 $X=180430 $Y=360750
X1462 963 1 966 953 2 ND2D1BWP7T $T=182960 364960 1 180 $X=180430 $Y=364725
X1463 954 1 310 973 2 ND2D1BWP7T $T=180720 396320 1 0 $X=180430 $Y=392110
X1464 939 1 313 963 2 ND2D1BWP7T $T=181280 372800 0 0 $X=180990 $Y=372565
X1465 947 1 302 932 2 ND2D1BWP7T $T=184640 372800 0 180 $X=182110 $Y=368590
X1466 980 1 315 961 2 ND2D1BWP7T $T=184640 388480 1 180 $X=182110 $Y=388245
X1467 969 1 925 313 2 ND2D1BWP7T $T=183520 372800 0 0 $X=183230 $Y=372565
X1468 963 1 971 961 2 ND2D1BWP7T $T=186320 388480 0 180 $X=183790 $Y=384270
X1469 964 1 318 978 2 ND2D1BWP7T $T=186880 388480 1 180 $X=184350 $Y=388245
X1470 961 1 319 932 2 ND2D1BWP7T $T=184640 396320 1 0 $X=184350 $Y=392110
X1471 941 1 322 264 2 ND2D1BWP7T $T=185760 404160 0 0 $X=185470 $Y=403925
X1472 963 1 291 947 2 ND2D1BWP7T $T=186320 372800 0 0 $X=186030 $Y=372565
X1473 972 1 316 948 2 ND2D1BWP7T $T=190240 388480 0 180 $X=187710 $Y=384270
X1474 963 1 326 948 2 ND2D1BWP7T $T=188560 372800 0 0 $X=188270 $Y=372565
X1475 964 1 332 319 2 ND2D1BWP7T $T=189680 396320 0 0 $X=189390 $Y=396085
X1476 972 1 306 947 2 ND2D1BWP7T $T=192480 388480 0 180 $X=189950 $Y=384270
X1477 985 1 329 994 2 ND2D1BWP7T $T=191920 372800 1 0 $X=191630 $Y=368590
X1478 973 1 264 972 2 ND2D1BWP7T $T=194720 388480 0 180 $X=192190 $Y=384270
X1479 998 1 340 1002 2 ND2D1BWP7T $T=194720 396320 0 0 $X=194430 $Y=396085
X1480 951 1 956 1002 2 ND2D1BWP7T $T=208160 380640 0 180 $X=205630 $Y=376430
X1481 998 1 345 993 2 ND2D1BWP7T $T=205920 396320 0 0 $X=205630 $Y=396085
X1482 1007 1 1000 1001 2 ND2D1BWP7T $T=210400 372800 0 180 $X=207870 $Y=368590
X1483 1002 1 1006 1007 2 ND2D1BWP7T $T=208160 372800 0 0 $X=207870 $Y=372565
X1484 1014 1 1003 1018 2 ND2D1BWP7T $T=219360 380640 1 0 $X=219070 $Y=376430
X1485 1018 1 1017 334 2 ND2D1BWP7T $T=226640 404160 0 0 $X=226350 $Y=403925
X1486 446 1 455 456 2 ND2D1BWP7T $T=296080 372800 1 0 $X=295790 $Y=368590
X1487 505 1 1085 456 2 ND2D1BWP7T $T=345920 380640 1 0 $X=345630 $Y=376430
X1488 160 1 834 805 2 803 863 OAI211D1BWP7T $T=86640 396320 1 0 $X=86350 $Y=392110
X1489 155 1 90 861 2 164 823 OAI211D1BWP7T $T=87760 412000 1 0 $X=87470 $Y=407790
X1490 160 1 834 805 2 879 863 OAI211D1BWP7T $T=94480 396320 1 0 $X=94190 $Y=392110
X1491 42 1 103 881 2 870 884 OAI211D1BWP7T $T=100640 372800 0 0 $X=100350 $Y=372565
X1492 896 1 830 897 2 205 898 OAI211D1BWP7T $T=111840 388480 1 0 $X=111550 $Y=384270
X1493 904 1 895 899 2 886 900 OAI211D1BWP7T $T=125280 364960 0 180 $X=121630 $Y=360750
X1494 868 1 182 211 2 902 900 OAI211D1BWP7T $T=121920 380640 1 0 $X=121630 $Y=376430
X1495 28 1 903 881 2 210 872 OAI211D1BWP7T $T=125840 372800 0 180 $X=122190 $Y=368590
X1496 895 1 904 899 2 213 900 OAI211D1BWP7T $T=128640 364960 0 180 $X=124990 $Y=360750
X1497 28 1 903 881 2 905 872 OAI211D1BWP7T $T=130880 364960 0 0 $X=130590 $Y=364725
X1498 316 1 328 245 2 325 992 OAI211D1BWP7T $T=188560 412000 0 0 $X=188270 $Y=411765
X1499 971 1 943 993 2 348 329 OAI211D1BWP7T $T=209280 404160 1 180 $X=205630 $Y=403925
X1500 915 1 359 334 2 1013 933 OAI211D1BWP7T $T=213200 404160 0 0 $X=212910 $Y=403925
X1501 275 1 943 1009 2 1015 1014 OAI211D1BWP7T $T=213760 388480 1 0 $X=213470 $Y=384270
X1502 943 1 366 1009 2 365 1017 OAI211D1BWP7T $T=217120 412000 1 0 $X=216830 $Y=407790
X1503 455 1 1068 1067 2 452 401 OAI211D1BWP7T $T=297760 380640 0 180 $X=294110 $Y=376430
X1504 1123 1 1119 1113 2 1110 542 OAI211D1BWP7T $T=367200 380640 1 180 $X=363550 $Y=380405
X1505 1146 1 1142 1141 2 1143 542 OAI211D1BWP7T $T=399680 388480 1 180 $X=396030 $Y=388245
X1506 1151 1 1149 582 2 1130 542 OAI211D1BWP7T $T=404160 380640 1 180 $X=400510 $Y=380405
X1507 828 2 808 49 38 1 50 NR4D2BWP7T $T=50800 388480 0 180 $X=37630 $Y=384270
X1508 808 2 807 792 794 1 826 NR4D2BWP7T $T=39040 380640 0 0 $X=38750 $Y=380405
X1509 38 2 819 56 802 1 59 NR4D2BWP7T $T=52480 396320 0 180 $X=39310 $Y=392110
X1510 128 2 847 841 792 1 99 NR4D2BWP7T $T=73200 396320 1 180 $X=60030 $Y=396085
X1511 838 2 889 794 810 1 830 NR4D2BWP7T $T=101200 396320 1 0 $X=100910 $Y=392110
X1512 912 2 913 233 928 1 238 NR4D2BWP7T $T=136480 412000 1 0 $X=136190 $Y=407790
X1513 55 2 7 817 1 NR2XD0BWP7T $T=44080 412000 1 0 $X=43790 $Y=407790
X1514 204 2 884 198 1 NR2XD0BWP7T $T=112960 357120 1 180 $X=110430 $Y=356885
X1515 18 1 790 791 788 793 2 ND4D1BWP7T $T=26720 380640 0 180 $X=22510 $Y=376430
X1516 68 1 42 821 59 62 2 ND4D1BWP7T $T=50240 364960 1 180 $X=46030 $Y=364725
X1517 69 1 790 47 822 813 2 ND4D1BWP7T $T=51360 372800 1 180 $X=47150 $Y=372565
X1518 834 1 81 825 74 832 2 ND4D1BWP7T $T=56960 388480 0 180 $X=52750 $Y=384270
X1519 79 1 826 17 845 120 2 ND4D1BWP7T $T=66480 372800 1 0 $X=66190 $Y=368590
X1520 121 1 117 825 833 852 2 ND4D1BWP7T $T=68160 364960 1 0 $X=67870 $Y=360750
X1521 42 1 152 855 822 147 2 ND4D1BWP7T $T=87200 372800 0 180 $X=82990 $Y=368590
X1522 107 1 169 862 94 866 2 ND4D1BWP7T $T=93360 388480 0 180 $X=89150 $Y=384270
X1523 921 1 917 915 229 912 2 ND4D1BWP7T $T=144320 404160 0 180 $X=140110 $Y=399950
X1524 922 1 261 258 926 251 2 ND4D1BWP7T $T=156640 404160 0 180 $X=152430 $Y=399950
X1525 261 1 262 936 254 913 2 ND4D1BWP7T $T=156640 412000 0 180 $X=152430 $Y=407790
X1526 270 1 302 969 966 970 2 ND4D1BWP7T $T=177360 372800 1 0 $X=177070 $Y=368590
X1527 941 1 310 316 981 323 2 ND4D1BWP7T $T=185200 412000 1 0 $X=184910 $Y=407790
X1528 306 1 981 971 976 988 2 ND4D1BWP7T $T=186320 404160 1 0 $X=186030 $Y=399950
X1529 971 1 955 1010 354 249 2 ND4D1BWP7T $T=209280 404160 0 0 $X=208990 $Y=403925
X1530 859 878 880 860 191 1 2 OAI31D1BWP7T $T=100640 364960 0 0 $X=100350 $Y=364725
X1531 852 905 212 891 215 1 2 OAI31D1BWP7T $T=124160 357120 0 0 $X=123870 $Y=356885
X1532 1001 999 997 990 937 1 2 OAI31D1BWP7T $T=196400 380640 1 180 $X=192190 $Y=380405
X1533 77 883 871 195 193 1 2 AOI31D0BWP7T $T=109040 412000 1 180 $X=105390 $Y=411765
X1534 103 1 104 74 2 836 ND3D0BWP7T $T=63120 372800 0 180 $X=60030 $Y=368590
X1535 864 1 166 826 2 860 ND3D0BWP7T $T=91120 364960 1 180 $X=88030 $Y=364725
X1536 865 1 167 834 2 878 ND3D0BWP7T $T=97280 380640 1 0 $X=96990 $Y=376430
X1537 300 1 286 971 2 968 ND3D0BWP7T $T=177920 388480 1 0 $X=177630 $Y=384270
X1538 93 1 2 817 827 837 95 NR4D0BWP7T $T=63120 404160 1 180 $X=59470 $Y=403925
X1539 101 1 2 129 159 151 846 NR4D0BWP7T $T=88880 364960 0 180 $X=85230 $Y=360750
X1540 129 1 2 165 820 864 163 NR4D0BWP7T $T=91120 357120 1 180 $X=87470 $Y=356885
X1541 839 1 2 819 199 896 859 NR4D0BWP7T $T=108480 388480 0 0 $X=108190 $Y=388245
X1542 253 1 2 249 231 250 242 NR4D0BWP7T $T=153280 412000 1 180 $X=149630 $Y=411765
X1543 927 1 2 968 314 978 931 NR4D0BWP7T $T=180720 388480 1 0 $X=180430 $Y=384270
X1544 1015 1 2 361 318 364 949 NR4D0BWP7T $T=218800 412000 1 180 $X=215150 $Y=411765
X1545 789 65 2 71 1 NR2D2BWP7T $T=47440 404160 0 0 $X=47150 $Y=403925
X1546 899 805 2 199 1 NR2D2BWP7T $T=122480 396320 1 0 $X=122190 $Y=392110
X1547 908 805 2 795 1 NR2D2BWP7T $T=130880 396320 1 180 $X=126670 $Y=396085
X1548 897 908 2 92 1 NR2D2BWP7T $T=136480 388480 1 180 $X=132270 $Y=388245
X1549 204 226 2 853 1 NR2D2BWP7T $T=142080 364960 1 180 $X=137870 $Y=364725
X1550 938 257 2 916 1 NR2D2BWP7T $T=157200 404160 1 180 $X=152990 $Y=403925
X1551 1006 993 2 972 1 NR2D2BWP7T $T=211520 357120 1 180 $X=207310 $Y=356885
X1552 1004 1009 2 297 1 NR2D2BWP7T $T=222720 404160 0 0 $X=222430 $Y=403925
X1553 916 982 319 264 2 1 336 AN4D1BWP7T $T=189680 404160 0 0 $X=189390 $Y=403925
X1554 975 1 2 976 BUFFD0BWP7T $T=179600 404160 1 0 $X=179310 $Y=399950
X1555 887 46 188 883 183 2 1 AOI31D1BWP7T $T=105680 412000 1 180 $X=101470 $Y=411765
X1556 920 73 890 227 842 2 1 AOI31D1BWP7T $T=143200 372800 0 180 $X=138990 $Y=368590
X1557 999 973 1010 1007 928 2 1 AOI31D1BWP7T $T=213200 388480 1 180 $X=208990 $Y=388245
X1558 42 1 39 36 31 798 2 ND4D0BWP7T $T=41280 357120 1 180 $X=37630 $Y=356885
X1559 47 1 28 44 41 804 2 ND4D0BWP7T $T=43520 372800 1 180 $X=39870 $Y=372565
X1560 18 1 68 824 825 66 2 ND4D0BWP7T $T=49120 372800 1 0 $X=48830 $Y=368590
X1561 94 1 788 44 834 835 2 ND4D0BWP7T $T=61440 388480 1 180 $X=57790 $Y=388245
X1562 124 1 825 850 86 132 2 ND4D0BWP7T $T=69840 357120 0 0 $X=69550 $Y=356885
X1563 201 1 892 873 41 891 2 ND4D0BWP7T $T=110160 357120 1 180 $X=106510 $Y=356885
X1564 893 1 169 895 834 208 2 ND4D0BWP7T $T=109040 372800 0 0 $X=108750 $Y=372565
X1565 280 1 283 284 957 958 2 ND4D0BWP7T $T=169520 404160 1 0 $X=169230 $Y=399950
X1566 315 1 302 294 316 320 2 ND4D0BWP7T $T=182400 412000 0 0 $X=182110 $Y=411765
X1567 310 1 945 279 306 986 2 ND4D0BWP7T $T=183520 396320 0 0 $X=183230 $Y=396085
X1568 844 1 890 2 893 196 IND3D1BWP7T $T=105680 372800 0 0 $X=105390 $Y=372565
X1569 154 148 93 2 1 NR2D1P5BWP7T $T=86640 412000 1 180 $X=82430 $Y=411765
X1570 19 127 884 2 1 NR2D1P5BWP7T $T=104000 396320 1 180 $X=99790 $Y=396085
X1571 55 183 206 2 1 NR2D1P5BWP7T $T=112960 412000 1 180 $X=108750 $Y=411765
X1572 934 276 956 2 1 NR2D1P5BWP7T $T=170640 396320 1 180 $X=166430 $Y=396085
X1573 1004 931 956 2 1 NR2D1P5BWP7T $T=199200 388480 1 180 $X=194990 $Y=388245
X1574 310 2 977 243 967 975 1 INR4D0BWP7T $T=186320 404160 0 180 $X=181550 $Y=399950
X1575 810 1 792 813 812 2 NR3D1BWP7T $T=42400 372800 1 0 $X=42110 $Y=368590
X1576 87 1 92 836 86 2 NR3D1BWP7T $T=60320 357120 1 180 $X=55550 $Y=356885
X1577 839 1 794 835 119 2 NR3D1BWP7T $T=61440 388480 0 0 $X=61150 $Y=388245
X1578 952 1 333 997 335 2 NR3D1BWP7T $T=195280 388480 1 180 $X=190510 $Y=388245
X1579 358 1 1011 988 360 2 NR3D1BWP7T $T=221040 404160 1 180 $X=216270 $Y=403925
X1580 838 1 873 152 876 824 2 IND4D0BWP7T $T=96720 388480 1 0 $X=96430 $Y=384270
X1581 273 1 945 270 266 264 2 IND4D0BWP7T $T=167840 412000 1 180 $X=163630 $Y=411765
X1582 257 1 288 283 960 291 2 IND4D0BWP7T $T=170640 372800 0 0 $X=170350 $Y=372565
X1583 128 1 854 138 135 43 2 IND4D1BWP7T $T=84400 357120 1 180 $X=79630 $Y=356885
X1584 832 2 829 63 16 1 58 NR4D3BWP7T $T=57520 388480 1 180 $X=41550 $Y=388245
X1585 879 882 153 190 868 1 2 INR4D1BWP7T $T=100640 388480 0 0 $X=100350 $Y=388245
X1586 842 889 214 216 28 1 2 INR4D1BWP7T $T=130320 372800 1 180 $X=123310 $Y=372565
X1587 184 173 851 903 104 1 2 INR4D1BWP7T $T=125840 380640 0 0 $X=125550 $Y=380405
X1588 231 923 927 917 240 1 2 INR4D1BWP7T $T=143760 396320 1 0 $X=143470 $Y=392110
X1589 983 321 935 2 1 INR2D2BWP7T $T=188560 357120 1 180 $X=183790 $Y=356885
X1590 3 2 789 1 12 NR2XD1BWP7T $T=21120 404160 0 0 $X=20830 $Y=403925
X1591 4 2 11 1 19 NR2XD1BWP7T $T=22800 357120 0 0 $X=22510 $Y=356885
X1592 799 2 802 1 805 NR2XD1BWP7T $T=26720 396320 1 0 $X=26430 $Y=392110
X1593 15 2 40 1 35 NR2XD1BWP7T $T=41840 412000 0 180 $X=37630 $Y=407790
X1594 15 2 811 1 800 NR2XD1BWP7T $T=39600 404160 1 0 $X=39310 $Y=399950
X1595 55 2 48 1 800 NR2XD1BWP7T $T=44640 404160 1 180 $X=40430 $Y=403925
X1596 15 2 65 1 823 NR2XD1BWP7T $T=46880 404160 1 0 $X=46590 $Y=399950
X1597 800 2 89 1 30 NR2XD1BWP7T $T=55280 404160 0 0 $X=54990 $Y=403925
X1598 6 2 93 1 35 NR2XD1BWP7T $T=57520 404160 1 0 $X=57230 $Y=399950
X1599 40 2 114 1 116 NR2XD1BWP7T $T=64240 404160 1 0 $X=63950 $Y=399950
X1600 823 2 116 1 30 NR2XD1BWP7T $T=72080 404160 0 180 $X=67870 $Y=399950
X1601 130 2 816 1 805 NR2XD1BWP7T $T=83840 396320 0 180 $X=79630 $Y=392110
X1602 811 2 139 1 26 NR2XD1BWP7T $T=83840 404160 0 180 $X=79630 $Y=399950
X1603 130 2 136 1 857 NR2XD1BWP7T $T=81040 396320 0 0 $X=80750 $Y=396085
X1604 823 2 162 1 6 NR2XD1BWP7T $T=85520 404160 1 0 $X=85230 $Y=399950
X1605 150 2 154 1 33 NR2XD1BWP7T $T=105680 404160 0 180 $X=101470 $Y=399950
X1606 35 2 203 1 150 NR2XD1BWP7T $T=113520 404160 0 180 $X=109310 $Y=399950
X1607 204 2 820 1 897 NR2XD1BWP7T $T=111280 364960 1 0 $X=110990 $Y=360750
X1608 884 2 21 1 899 NR2XD1BWP7T $T=111280 364960 0 0 $X=110990 $Y=364725
X1609 899 2 814 1 857 NR2XD1BWP7T $T=115200 396320 1 180 $X=110990 $Y=396085
X1610 202 2 78 1 887 NR2XD1BWP7T $T=115200 412000 0 180 $X=110990 $Y=407790
X1611 897 2 841 1 863 NR2XD1BWP7T $T=126400 388480 1 180 $X=122190 $Y=388245
X1612 906 2 877 1 871 NR2XD1BWP7T $T=138160 404160 0 180 $X=133950 $Y=399950
X1613 235 2 237 1 929 NR2XD1BWP7T $T=146560 388480 0 0 $X=146270 $Y=388245
X1614 235 2 231 1 239 NR2XD1BWP7T $T=147680 404160 1 0 $X=147390 $Y=399950
X1615 226 2 848 1 236 NR2XD1BWP7T $T=153280 372800 0 180 $X=149070 $Y=368590
X1616 934 2 244 1 239 NR2XD1BWP7T $T=153280 404160 1 180 $X=149070 $Y=403925
X1617 930 2 252 1 256 NR2XD1BWP7T $T=151040 380640 1 0 $X=150750 $Y=376430
X1618 263 2 257 1 930 NR2XD1BWP7T $T=156640 372800 1 180 $X=152430 $Y=372565
X1619 946 2 943 1 252 NR2XD1BWP7T $T=167840 372800 1 180 $X=163630 $Y=372565
X1620 321 2 953 1 983 NR2XD1BWP7T $T=193040 357120 1 180 $X=188830 $Y=356885
X1621 990 2 337 1 245 NR2XD1BWP7T $T=191920 412000 0 0 $X=191630 $Y=411765
X1622 339 2 985 1 983 NR2XD1BWP7T $T=197520 357120 1 180 $X=193310 $Y=356885
X1623 929 2 342 1 990 NR2XD1BWP7T $T=198640 388480 0 180 $X=194430 $Y=384270
X1624 1000 2 944 1 999 NR2XD1BWP7T $T=199200 372800 0 180 $X=194990 $Y=368590
X1625 990 2 343 1 239 NR2XD1BWP7T $T=195280 412000 1 0 $X=194990 $Y=407790
X1626 345 2 954 1 1002 NR2XD1BWP7T $T=205920 396320 1 0 $X=205630 $Y=392110
X1627 345 2 980 1 1001 NR2XD1BWP7T $T=206480 380640 0 0 $X=206190 $Y=380405
X1628 1007 2 951 1 993 NR2XD1BWP7T $T=214320 372800 1 180 $X=210110 $Y=372565
X1629 1004 2 358 1 245 NR2XD1BWP7T $T=216560 404160 0 180 $X=212350 $Y=399950
X1630 1003 2 965 1 334 NR2XD1BWP7T $T=218240 372800 1 180 $X=214030 $Y=372565
X1631 1009 2 362 1 256 NR2XD1BWP7T $T=220480 396320 0 180 $X=216270 $Y=392110
X1632 810 1 129 833 2 IND2D1BWP7T $T=73200 364960 1 180 $X=70110 $Y=364725
X1633 177 1 869 61 2 IND2D1BWP7T $T=96720 357120 1 180 $X=93630 $Y=356885
X1634 794 1 200 895 2 IND2D1BWP7T $T=108480 364960 0 0 $X=108190 $Y=364725
X1635 92 1 101 904 2 IND2D1BWP7T $T=131440 380640 0 180 $X=128350 $Y=376430
X1636 923 1 952 286 2 IND2D1BWP7T $T=169520 380640 1 0 $X=169230 $Y=376430
X1637 925 1 1011 943 2 IND2D1BWP7T $T=209840 404160 1 0 $X=209550 $Y=399950
X1638 1005 1011 273 362 2 1 367 OR4XD1BWP7T $T=214880 396320 0 0 $X=214590 $Y=396085
X1639 28 1 903 881 2 872 220 OAI211D0BWP7T $T=126960 364960 0 0 $X=126670 $Y=364725
X1640 790 1 788 19 23 20 2 OAI211D2BWP7T $T=22240 388480 0 0 $X=21950 $Y=388245
X1641 969 1 981 321 331 987 2 OAI211D2BWP7T $T=185200 372800 1 0 $X=184910 $Y=368590
X1642 981 1 356 1014 353 239 2 OAI211D2BWP7T $T=213760 380640 0 0 $X=213470 $Y=380405
X1643 1085 1 1089 401 1020 1079 2 OAI211D2BWP7T $T=322400 380640 1 180 $X=315950 $Y=380405
X1644 1085 1 1118 401 535 1112 2 OAI211D2BWP7T $T=363280 388480 1 180 $X=356830 $Y=388245
X1645 815 877 811 789 1 2 185 AO211D0BWP7T $T=98400 412000 1 0 $X=98110 $Y=407790
X1646 849 73 882 875 1 2 874 AO211D0BWP7T $T=106800 372800 0 180 $X=102590 $Y=368590
X1647 225 849 223 909 1 2 222 AO211D0BWP7T $T=135920 357120 1 180 $X=131710 $Y=356885
X1648 961 951 925 960 1 2 984 AO211D0BWP7T $T=184640 380640 1 0 $X=184350 $Y=376430
X1649 985 954 318 986 1 2 995 AO211D0BWP7T $T=190240 396320 1 0 $X=189950 $Y=392110
X1650 122 2 126 115 843 9 1 AOI211D2BWP7T $T=70960 380640 0 180 $X=64510 $Y=376430
X1651 322 2 324 338 996 993 1 AOI211D2BWP7T $T=189120 412000 1 0 $X=188830 $Y=407790
X1652 15 2 10 7 1 NR2D3BWP7T $T=27280 412000 1 180 $X=21950 $Y=411765
X1653 12 2 29 30 1 NR2D3BWP7T $T=25040 404160 0 0 $X=24750 $Y=403925
X1654 6 2 26 12 1 NR2D3BWP7T $T=31200 404160 0 180 $X=25870 $Y=399950
X1655 800 2 113 45 1 NR2D3BWP7T $T=69840 412000 0 180 $X=64510 $Y=407790
X1656 871 2 34 202 1 NR2D3BWP7T $T=106240 404160 0 0 $X=105950 $Y=403925
X1657 897 2 122 19 1 NR2D3BWP7T $T=115200 380640 0 180 $X=109870 $Y=376430
X1658 897 2 810 910 1 NR2D3BWP7T $T=128080 396320 1 0 $X=127790 $Y=392110
X1659 861 2 224 871 1 NR2D3BWP7T $T=131440 412000 1 0 $X=131150 $Y=407790
X1660 20 2 27 226 1 NR2D3BWP7T $T=144320 380640 1 180 $X=138990 $Y=380405
X1661 918 2 5 226 1 NR2D3BWP7T $T=148240 380640 0 180 $X=142910 $Y=376430
X1662 881 2 809 234 1 NR2D3BWP7T $T=151600 364960 1 180 $X=146270 $Y=364725
X1663 235 2 248 933 1 NR2D3BWP7T $T=148240 396320 0 0 $X=147950 $Y=396085
X1664 1003 2 947 994 1 NR2D3BWP7T $T=198080 372800 1 180 $X=192750 $Y=372565
X1665 1004 2 304 933 1 NR2D3BWP7T $T=199200 396320 0 180 $X=193870 $Y=392110
X1666 1006 2 963 999 1 NR2D3BWP7T $T=208160 364960 0 0 $X=207870 $Y=364725
X1667 992 2 973 1018 1 NR2D3BWP7T $T=219360 388480 1 0 $X=219070 $Y=384270
X1668 934 2 273 1009 1 NR2D3BWP7T $T=222160 396320 1 0 $X=221870 $Y=392110
X1669 73 848 1 2 898 221 884 MOAI22D0BWP7T $T=134240 372800 0 180 $X=130030 $Y=368590
X1670 980 965 1 2 305 AN2D1BWP7T $T=209840 396320 1 0 $X=209550 $Y=392110
X1671 8 22 797 1 2 ND2D2BWP7T $T=25600 372800 0 0 $X=25310 $Y=372565
X1672 27 57 797 1 2 ND2D2BWP7T $T=43520 380640 1 0 $X=43230 $Y=376430
X1673 871 6 178 1 2 ND2D2BWP7T $T=97840 404160 0 180 $X=93630 $Y=399950
X1674 883 45 877 1 2 ND2D2BWP7T $T=106240 404160 1 180 $X=102030 $Y=403925
X1675 207 35 85 1 2 ND2D2BWP7T $T=115200 404160 1 180 $X=110990 $Y=403925
X1676 85 800 217 1 2 ND2D2BWP7T $T=128080 412000 1 180 $X=123870 $Y=411765
X1677 901 150 907 1 2 ND2D2BWP7T $T=125840 404160 1 0 $X=125550 $Y=399950
X1678 877 219 907 1 2 ND2D2BWP7T $T=130880 404160 1 180 $X=126670 $Y=403925
X1679 848 884 920 1 2 ND2D2BWP7T $T=143200 372800 1 0 $X=142910 $Y=368590
X1680 980 279 947 1 2 ND2D2BWP7T $T=186880 388480 0 0 $X=186590 $Y=388245
X1681 1001 245 951 1 2 ND2D2BWP7T $T=213200 380640 0 180 $X=208990 $Y=376430
X1682 1016 256 983 1 2 ND2D2BWP7T $T=222160 372800 1 180 $X=217950 $Y=372565
X1683 816 1 2 126 149 858 NR3D0BWP7T $T=83280 388480 0 0 $X=82990 $Y=388245
X1684 63 1 2 820 875 181 NR3D0BWP7T $T=97840 357120 0 0 $X=97550 $Y=356885
X1685 1003 263 1 929 1005 2 AOI21D1BWP7T $T=199200 380640 0 180 $X=195550 $Y=376430
X1686 529 1098 1 1105 1103 2 AOI21D1BWP7T $T=352640 404160 1 180 $X=348990 $Y=403925
X1687 503 1137 1 576 1120 2 AOI21D1BWP7T $T=389040 388480 1 0 $X=388750 $Y=384270
X1688 596 1145 1 1158 1155 2 AOI21D1BWP7T $T=424320 357120 1 180 $X=420670 $Y=356885
X1689 80 865 177 169 2 1 ND3D2BWP7T $T=92240 380640 0 0 $X=91950 $Y=380405
X1690 259 241 910 230 2 1 ND3D2BWP7T $T=157200 357120 1 180 $X=151870 $Y=356885
X1691 858 44 824 121 153 1 2 ND4D2BWP7T $T=87200 388480 0 180 $X=79630 $Y=384270
X1692 57 167 862 68 171 1 2 ND4D2BWP7T $T=88880 372800 0 0 $X=88590 $Y=372565
X1693 80 1 57 830 2 828 ND3D1BWP7T $T=55280 380640 1 180 $X=51630 $Y=380405
X1694 88 1 90 71 2 84 ND3D1BWP7T $T=56400 412000 0 0 $X=56110 $Y=411765
X1695 865 1 124 137 2 128 ND3D1BWP7T $T=90560 372800 0 180 $X=86910 $Y=368590
X1696 922 1 919 916 2 228 ND3D1BWP7T $T=144320 412000 1 180 $X=140670 $Y=411765
X1697 67 2 63 818 1 821 9 AOI211D1BWP7T $T=50800 364960 0 180 $X=47150 $Y=360750
X1698 793 2 829 853 1 854 142 AOI211D1BWP7T $T=79920 372800 1 0 $X=79630 $Y=368590
X1699 875 2 198 894 1 892 831 AOI211D1BWP7T $T=107920 364960 1 0 $X=107630 $Y=360750
X1700 327 2 952 985 1 982 932 AOI211D1BWP7T $T=190240 396320 0 180 $X=186590 $Y=392110
X1701 304 2 967 998 1 341 996 AOI211D1BWP7T $T=193600 404160 1 0 $X=193310 $Y=399950
X1702 1080 2 1078 1049 1 1068 487 AOI211D1BWP7T $T=317360 372800 1 180 $X=313710 $Y=372565
X1703 1115 2 541 1116 1 1119 391 AOI211D1BWP7T $T=359360 380640 1 0 $X=359070 $Y=376430
X1704 547 2 541 1107 1 1126 391 AOI211D1BWP7T $T=377280 364960 1 0 $X=376990 $Y=360750
X1705 1 2 ICV_17 $T=52480 396320 1 0 $X=52190 $Y=392110
X1706 1 2 ICV_17 $T=56960 412000 1 0 $X=56670 $Y=407790
X1707 1 2 ICV_17 $T=119120 412000 0 0 $X=118830 $Y=411765
X1708 1 2 ICV_17 $T=131440 380640 1 0 $X=131150 $Y=376430
X1709 1 2 ICV_17 $T=133120 388480 1 0 $X=132830 $Y=384270
X1710 1 2 ICV_17 $T=312320 404160 0 0 $X=312030 $Y=403925
X1711 1 2 ICV_17 $T=313440 357120 0 0 $X=313150 $Y=356885
X1712 1 2 ICV_17 $T=313440 396320 0 0 $X=313150 $Y=396085
X1713 1 2 ICV_17 $T=344800 388480 0 0 $X=344510 $Y=388245
X1714 1 2 ICV_17 $T=347600 364960 0 0 $X=347310 $Y=364725
X1715 1 2 ICV_17 $T=352080 388480 0 0 $X=351790 $Y=388245
X1716 1 2 ICV_17 $T=358800 380640 0 0 $X=358510 $Y=380405
X1717 1 2 ICV_17 $T=359920 396320 0 0 $X=359630 $Y=396085
X1718 1 2 ICV_17 $T=383440 380640 1 0 $X=383150 $Y=376430
X1719 1 2 ICV_17 $T=422080 364960 1 0 $X=421790 $Y=360750
X1720 1 2 ICV_17 $T=423200 396320 1 0 $X=422910 $Y=392110
X1721 1 2 ICV_17 $T=463520 388480 1 0 $X=463230 $Y=384270
X1739 33 12 2 1 CKBD2BWP7T $T=31200 396320 1 180 $X=27550 $Y=396085
X1740 651 462 2 1 CKBD2BWP7T $T=464640 372800 0 180 $X=460990 $Y=368590
X1741 1172 643 641 1174 544 1 2 1175 AO221D0BWP7T $T=459040 404160 1 0 $X=458750 $Y=399950
X1742 1 2 ICV_19 $T=27840 364960 1 0 $X=27550 $Y=360750
X1743 1 2 ICV_19 $T=153840 364960 1 0 $X=153550 $Y=360750
X1744 1 2 ICV_19 $T=182960 364960 1 0 $X=182670 $Y=360750
X1745 1 2 ICV_19 $T=237840 364960 1 0 $X=237550 $Y=360750
X1746 1 2 ICV_19 $T=237840 396320 0 0 $X=237550 $Y=396085
X1747 1 2 ICV_19 $T=237840 404160 1 0 $X=237550 $Y=399950
X1748 1 2 ICV_19 $T=237840 404160 0 0 $X=237550 $Y=403925
X1749 1 2 ICV_19 $T=262480 396320 0 0 $X=262190 $Y=396085
X1750 1 2 ICV_19 $T=272560 412000 1 0 $X=272270 $Y=407790
X1751 1 2 ICV_19 $T=304480 357120 0 0 $X=304190 $Y=356885
X1752 1 2 ICV_19 $T=321840 372800 1 0 $X=321550 $Y=368590
X1753 1 2 ICV_19 $T=321840 412000 1 0 $X=321550 $Y=407790
X1754 1 2 ICV_19 $T=363840 412000 1 0 $X=363550 $Y=407790
X1755 1 2 ICV_19 $T=392400 372800 1 0 $X=392110 $Y=368590
X1756 1 2 ICV_19 $T=438320 364960 1 0 $X=438030 $Y=360750
X1757 1 2 ICV_19 $T=447840 380640 1 0 $X=447550 $Y=376430
X1758 1 2 ICV_19 $T=447840 388480 0 0 $X=447550 $Y=388245
X1759 1 2 ICV_19 $T=455120 372800 1 0 $X=454830 $Y=368590
X1778 1 2 ICV_21 $T=26720 372800 1 0 $X=26430 $Y=368590
X1779 1 2 ICV_21 $T=47440 380640 1 0 $X=47150 $Y=376430
X1780 1 2 ICV_21 $T=104000 412000 1 0 $X=103710 $Y=407790
X1781 1 2 ICV_21 $T=236720 372800 0 0 $X=236430 $Y=372565
X1782 1 2 ICV_21 $T=273120 412000 0 0 $X=272830 $Y=411765
X1783 1 2 ICV_21 $T=278720 388480 0 0 $X=278430 $Y=388245
X1784 1 2 ICV_21 $T=278720 404160 1 0 $X=278430 $Y=399950
X1785 1 2 ICV_21 $T=291600 364960 0 0 $X=291310 $Y=364725
X1786 1 2 ICV_21 $T=304480 412000 0 0 $X=304190 $Y=411765
X1787 1 2 ICV_21 $T=306720 372800 0 0 $X=306430 $Y=372565
X1788 1 2 ICV_21 $T=329120 380640 1 0 $X=328830 $Y=376430
X1789 1 2 ICV_21 $T=380640 364960 1 0 $X=380350 $Y=360750
X1790 1 2 ICV_21 $T=381760 388480 1 0 $X=381470 $Y=384270
X1791 1 2 ICV_21 $T=385120 372800 0 0 $X=384830 $Y=372565
X1792 1 2 ICV_21 $T=436640 404160 1 0 $X=436350 $Y=399950
X1793 1 2 ICV_21 $T=446720 388480 1 0 $X=446430 $Y=384270
X1794 1 2 ICV_21 $T=446720 404160 1 0 $X=446430 $Y=399950
X1799 436 1165 532 599 2 1 1161 DFCND1BWP7T $T=437760 372800 1 180 $X=424590 $Y=372565
X1800 400 394 906 1 2 XNR2D2BWP7T $T=239520 388480 0 180 $X=232510 $Y=384270
X1801 490 478 999 1 2 XNR2D2BWP7T $T=316240 364960 0 180 $X=309230 $Y=360750
X1802 508 502 1002 1 2 XNR2D2BWP7T $T=325200 357120 1 180 $X=318190 $Y=356885
X1803 538 1110 533 1 2 XNR2D2BWP7T $T=361600 364960 0 180 $X=354590 $Y=360750
X1804 606 1143 998 1 2 XNR2D2BWP7T $T=427680 404160 0 180 $X=420670 $Y=399950
X1805 789 1 2 827 34 82 85 AOI211XD0BWP7T $T=53600 412000 1 0 $X=53310 $Y=407790
X1806 840 1 2 846 848 161 9 AOI211XD0BWP7T $T=83280 364960 0 0 $X=82990 $Y=364725
X1807 162 1 2 113 815 174 178 AOI211XD0BWP7T $T=92240 412000 1 0 $X=91950 $Y=407790
X1808 184 1 2 802 885 888 806 AOI211XD0BWP7T $T=101760 380640 1 0 $X=101470 $Y=376430
X1809 131 1 2 886 831 194 885 AOI211XD0BWP7T $T=104000 364960 1 0 $X=103710 $Y=360750
X1810 1147 1 2 588 1138 1156 391 AOI211XD0BWP7T $T=400800 380640 1 0 $X=400510 $Y=376430
X1811 1155 1 2 593 583 1149 391 AOI211XD0BWP7T $T=409200 357120 1 180 $X=405550 $Y=356885
X1812 1163 1 2 588 1159 1142 391 AOI211XD0BWP7T $T=422640 388480 1 180 $X=418990 $Y=388245
X1813 372 1040 380 408 406 1 2 DFCND2BWP7T $T=266400 364960 0 180 $X=251550 $Y=360750
X1814 372 1032 380 1176 412 1 2 DFCND2BWP7T $T=252960 357120 0 0 $X=252670 $Y=356885
X1815 372 1042 380 424 1044 1 2 DFCND2BWP7T $T=261360 364960 0 0 $X=261070 $Y=364725
X1816 436 1070 380 1052 1177 1 2 DFCND2BWP7T $T=310640 388480 0 180 $X=295790 $Y=384270
X1817 436 608 532 594 1152 1 2 DFCND2BWP7T $T=431040 372800 0 180 $X=416190 $Y=368590
X1818 849 1 822 9 797 2 OAI21D2BWP7T $T=72640 388480 0 180 $X=67310 $Y=384270
X1819 895 1 159 130 897 2 OAI21D2BWP7T $T=134240 364960 1 0 $X=133950 $Y=360750
X1820 167 1 184 884 910 2 OAI21D2BWP7T $T=134240 372800 1 0 $X=133950 $Y=368590
X1821 1128 1 553 559 1132 2 OAI21D2BWP7T $T=376720 357120 0 0 $X=376430 $Y=356885
X1822 598 1 595 559 1157 2 OAI21D2BWP7T $T=420960 357120 1 180 $X=415630 $Y=356885
X1823 1076 404 1 485 1074 2 IOA21D1BWP7T $T=314560 372800 0 180 $X=310910 $Y=368590
X1824 1153 558 1 1035 590 2 IOA21D1BWP7T $T=406400 404160 1 180 $X=402750 $Y=403925
X1825 1148 542 1 587 2 1147 1144 OAI22D1BWP7T $T=402480 372800 0 180 $X=398270 $Y=368590
X1826 567 1 2 1129 DEL1BWP7T $T=385120 388480 1 180 $X=379230 $Y=388245
X1827 524 1081 1065 1121 544 1 2 1122 AO221D1BWP7T $T=361600 404160 0 0 $X=361310 $Y=403925
X1828 530 529 1063 543 544 1 2 546 AO221D1BWP7T $T=361600 412000 0 0 $X=361310 $Y=411765
X1829 527 539 1072 1127 544 1 2 1134 AO221D1BWP7T $T=378960 412000 1 0 $X=378670 $Y=407790
X1830 372 374 380 1178 2 1 392 DFCND0BWP7T $T=222160 357120 0 0 $X=221870 $Y=356885
X1831 372 1048 380 1057 2 1 1059 DFCND0BWP7T $T=267520 372800 0 0 $X=267230 $Y=372565
X1832 372 1051 380 1055 2 1 1179 DFCND0BWP7T $T=268640 380640 0 0 $X=268350 $Y=380405
X1833 436 1077 494 1086 2 1 1083 DFCND0BWP7T $T=311760 396320 1 0 $X=311470 $Y=392110
X1834 436 1091 494 1094 2 1 1092 DFCND0BWP7T $T=347040 396320 0 180 $X=333870 $Y=392110
X1835 436 1104 494 1108 2 1 1109 DFCND0BWP7T $T=342000 404160 1 0 $X=341710 $Y=399950
X1836 436 1106 532 1099 2 1 1111 DFCND0BWP7T $T=349280 372800 1 0 $X=348990 $Y=368590
X1837 436 1102 532 1180 2 1 1100 DFCND0BWP7T $T=352640 364960 0 0 $X=352350 $Y=364725
X1838 444 409 435 1060 431 424 2 1054 1 OA222D0BWP7T $T=283200 364960 1 180 $X=276750 $Y=364725
X1839 525 493 435 1086 433 1094 2 1090 1 OA222D0BWP7T $T=340880 388480 0 180 $X=334430 $Y=384270
X1840 511 409 435 1094 433 1060 2 1101 1 OA222D0BWP7T $T=335280 380640 0 0 $X=334990 $Y=380405
X1841 512 409 435 1099 433 1086 2 1082 1 OA222D0BWP7T $T=342560 380640 0 180 $X=336110 $Y=376430
X1842 523 409 435 1056 433 1099 2 1097 1 OA222D0BWP7T $T=344800 372800 0 180 $X=338350 $Y=368590
X1843 125 2 141 1 157 145 85 AOI211XD1BWP7T $T=81600 404160 0 0 $X=81310 $Y=403925
X1844 1096 2 1103 1 1089 487 1098 AOI211XD1BWP7T $T=343120 396320 1 180 $X=336110 $Y=396085
X1845 34 30 1 2 INVD2P5BWP7T $T=31200 412000 0 180 $X=28110 $Y=407790
X1846 481 443 1 2 INVD2P5BWP7T $T=310640 357120 0 0 $X=310350 $Y=356885
X1847 461 464 1 2 INVD6BWP7T $T=298880 364960 0 0 $X=298590 $Y=364725
X1848 409 443 1 435 1056 431 429 2 1048 OAI222D2BWP7T $T=282080 357120 1 180 $X=271710 $Y=356885
X1849 409 1063 1 435 408 433 1052 2 1040 OAI222D2BWP7T $T=282640 380640 0 180 $X=272270 $Y=376430
X1850 409 1065 1 435 434 433 432 2 1051 OAI222D2BWP7T $T=283200 388480 0 180 $X=272830 $Y=384270
X1851 409 1072 1 435 1052 433 434 2 1070 OAI222D2BWP7T $T=302800 380640 1 180 $X=292430 $Y=380405
X1852 404 1 2 409 INVD5BWP7T $T=251840 372800 1 0 $X=251550 $Y=368590
X1853 373 370 207 1 2 XOR2D2BWP7T $T=225520 372800 0 180 $X=218510 $Y=368590
X1854 900 2 1 226 818 NR2D2P5BWP7T $T=143760 396320 0 180 $X=138430 $Y=392110
X1855 956 2 1 256 255 NR2D2P5BWP7T $T=175120 388480 0 180 $X=169790 $Y=384270
X1856 993 2 1 1000 932 NR2D2P5BWP7T $T=198640 364960 0 180 $X=193310 $Y=360750
X1857 339 994 956 991 326 1 2 OAI31D0BWP7T $T=195840 380640 0 180 $X=192190 $Y=376430
X1858 5 9 794 2 1 CKAN2D2BWP7T $T=21680 372800 0 0 $X=21390 $Y=372565
X1859 334 985 939 2 1 CKAN2D2BWP7T $T=193040 364960 0 180 $X=188830 $Y=360750
X1860 932 953 1 2 314 CKAN2D1BWP7T $T=182960 364960 0 0 $X=182670 $Y=364725
X1861 973 263 1 2 CKND4BWP7T $T=182400 380640 0 180 $X=178190 $Y=376430
X1862 957 926 286 293 2 1 962 AN4D0BWP7T $T=172320 404160 0 0 $X=172030 $Y=403925
X1863 970 2 952 946 292 1 NR3D2BWP7T $T=175680 364960 1 180 $X=165310 $Y=364725
X1864 259 863 204 1 2 OR2D2BWP7T $T=155520 364960 1 180 $X=151310 $Y=364725
X1865 245 256 931 229 2 1 IAO21D2BWP7T $T=155520 388480 1 180 $X=150190 $Y=388245
X1866 5 28 797 1 2 ND2D1P5BWP7T $T=31200 380640 0 180 $X=26990 $Y=376430
X1867 883 55 901 1 2 ND2D1P5BWP7T $T=121920 404160 1 0 $X=121630 $Y=399950
X1868 226 805 911 1 2 ND2D1P5BWP7T $T=138720 396320 1 180 $X=134510 $Y=396085
X1869 840 822 118 144 1 2 829 IIND4D1BWP7T $T=86080 372800 1 180 $X=80190 $Y=372565
X1870 36 41 810 1 2 INR2XD1BWP7T $T=38480 364960 1 0 $X=38190 $Y=360750
X1871 134 140 789 1 2 INR2XD1BWP7T $T=79920 412000 1 0 $X=79630 $Y=407790
X1872 805 91 1 2 INVD1P5BWP7T $T=59760 396320 0 180 $X=57230 $Y=392110
X1873 100 2 792 843 1 118 797 AOI211XD2BWP7T $T=57520 380640 0 0 $X=57230 $Y=380405
X1874 4 2 1 792 799 NR2XD2BWP7T $T=21120 364960 1 0 $X=20830 $Y=360750
X1875 6 2 1 13 800 NR2XD2BWP7T $T=21120 396320 0 0 $X=20830 $Y=396085
.ENDS
***************************************
.SUBCKT CKND6BWP7T I ZN VSS VDD
** N=4 EP=4 IP=0 FDC=11
M0 ZN I VSS VSS N L=1.8e-07 W=7.9e-07 $X=2080 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=7.9e-07 $X=2800 $Y=345 $D=0
M2 ZN I VSS VSS N L=1.8e-07 W=7.9e-07 $X=3520 $Y=345 $D=0
M3 VSS I ZN VSS N L=1.8e-07 W=7.9e-07 $X=4240 $Y=345 $D=0
M4 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=640 $Y=2205 $D=16
M5 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1360 $Y=2205 $D=16
M6 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=2080 $Y=2205 $D=16
M7 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=2800 $Y=2205 $D=16
M8 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=3520 $Y=2205 $D=16
M9 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=4240 $Y=2205 $D=16
D10 VSS I DN AREA=2.037e-13 PJ=1.81e-06 $X=140 $Y=860 $D=32
.ENDS
***************************************
.SUBCKT OAI221D2BWP7T C VSS B1 B2 ZN A2 VDD A1
** N=14 EP=8 IP=0 FDC=20
M0 VSS C 9 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 9 C VSS VSS N L=1.8e-07 W=1e-06 $X=1420 $Y=345 $D=0
M2 10 B2 9 VSS N L=1.8e-07 W=1e-06 $X=2140 $Y=345 $D=0
M3 9 B1 10 VSS N L=1.8e-07 W=1e-06 $X=2860 $Y=345 $D=0
M4 10 B1 9 VSS N L=1.8e-07 W=1e-06 $X=3580 $Y=345 $D=0
M5 9 B2 10 VSS N L=1.8e-07 W=1e-06 $X=4300 $Y=345 $D=0
M6 10 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=5800 $Y=345 $D=0
M7 ZN A2 10 VSS N L=1.8e-07 W=1e-06 $X=6520 $Y=345 $D=0
M8 10 A2 ZN VSS N L=1.8e-07 W=1e-06 $X=7280 $Y=345 $D=0
M9 ZN A1 10 VSS N L=1.8e-07 W=1e-06 $X=8040 $Y=345 $D=0
M10 VDD C ZN VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M11 ZN C VDD VDD P L=1.8e-07 W=1.37e-06 $X=1420 $Y=2205 $D=16
M12 11 B2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2180 $Y=2205 $D=16
M13 VDD B1 11 VDD P L=1.8e-07 W=1.37e-06 $X=2860 $Y=2205 $D=16
M14 12 B1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3660 $Y=2205 $D=16
M15 ZN B2 12 VDD P L=1.8e-07 W=1.37e-06 $X=4260 $Y=2205 $D=16
M16 13 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=5900 $Y=2205 $D=16
M17 VDD A2 13 VDD P L=1.8e-07 W=1.37e-06 $X=6520 $Y=2205 $D=16
M18 14 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=7320 $Y=2205 $D=16
M19 ZN A1 14 VDD P L=1.8e-07 W=1.37e-06 $X=7930 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_23 1 2
** N=2 EP=2 IP=4 FDC=10
X0 1 2 DCAP4BWP7T $T=4480 0 0 0 $X=4190 $Y=-235
X1 1 2 DCAP8BWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT INVD8BWP7T I ZN VSS VDD
** N=4 EP=4 IP=0 FDC=16
M0 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=715 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=1435 $Y=345 $D=0
M2 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=2175 $Y=345 $D=0
M3 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=2895 $Y=345 $D=0
M4 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=3635 $Y=345 $D=0
M5 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=4355 $Y=345 $D=0
M6 ZN I VSS VSS N L=1.8e-07 W=1e-06 $X=5095 $Y=345 $D=0
M7 VSS I ZN VSS N L=1.8e-07 W=1e-06 $X=5815 $Y=345 $D=0
M8 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=715 $Y=2205 $D=16
M9 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1435 $Y=2205 $D=16
M10 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=2175 $Y=2205 $D=16
M11 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=2895 $Y=2205 $D=16
M12 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=3635 $Y=2205 $D=16
M13 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=4355 $Y=2205 $D=16
M14 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=5095 $Y=2205 $D=16
M15 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=5815 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AO22D0BWP7T B2 A1 A2 B1 VSS VDD Z
** N=11 EP=7 IP=0 FDC=10
M0 10 B2 VSS VSS N L=1.8e-07 W=5e-07 $X=620 $Y=460 $D=0
M1 8 B1 10 VSS N L=1.8e-07 W=5e-07 $X=1115 $Y=460 $D=0
M2 11 A1 8 VSS N L=1.8e-07 W=5e-07 $X=1915 $Y=460 $D=0
M3 VSS A2 11 VSS N L=1.8e-07 W=5e-07 $X=2475 $Y=460 $D=0
M4 Z 8 VSS VSS N L=1.8e-07 W=5e-07 $X=3675 $Y=460 $D=0
M5 9 B2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2670 $D=16
M6 8 A1 9 VDD P L=1.8e-07 W=6.85e-07 $X=1415 $Y=2670 $D=16
M7 9 A2 8 VDD P L=1.8e-07 W=6.85e-07 $X=2235 $Y=2670 $D=16
M8 VDD B1 9 VDD P L=1.8e-07 W=6.85e-07 $X=2955 $Y=2670 $D=16
M9 Z 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=3675 $Y=2670 $D=16
.ENDS
***************************************
.SUBCKT CKND10BWP7T I VDD ZN VSS
** N=4 EP=4 IP=0 FDC=18
M0 ZN I VSS VSS N L=1.8e-07 W=6.55e-07 $X=1340 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=6.55e-07 $X=2060 $Y=345 $D=0
M2 ZN I VSS VSS N L=1.8e-07 W=6.55e-07 $X=2780 $Y=345 $D=0
M3 VSS I ZN VSS N L=1.8e-07 W=6.55e-07 $X=3500 $Y=345 $D=0
M4 ZN I VSS VSS N L=1.8e-07 W=6.55e-07 $X=4220 $Y=345 $D=0
M5 VSS I ZN VSS N L=1.8e-07 W=6.55e-07 $X=4940 $Y=345 $D=0
M6 ZN I VSS VSS N L=1.8e-07 W=6.55e-07 $X=5660 $Y=345 $D=0
M7 VSS I ZN VSS N L=1.8e-07 W=6.55e-07 $X=6380 $Y=345 $D=0
M8 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M9 VDD I ZN VDD P L=1.8e-07 W=1.565e-06 $X=1340 $Y=2010 $D=16
M10 ZN I VDD VDD P L=1.8e-07 W=1.565e-06 $X=2060 $Y=2010 $D=16
M11 VDD I ZN VDD P L=1.8e-07 W=1.565e-06 $X=2780 $Y=2010 $D=16
M12 ZN I VDD VDD P L=1.8e-07 W=1.565e-06 $X=3500 $Y=2010 $D=16
M13 VDD I ZN VDD P L=1.8e-07 W=1.565e-06 $X=4220 $Y=2010 $D=16
M14 ZN I VDD VDD P L=1.8e-07 W=1.565e-06 $X=4940 $Y=2010 $D=16
M15 VDD I ZN VDD P L=1.8e-07 W=1.565e-06 $X=5660 $Y=2010 $D=16
M16 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=6380 $Y=2205 $D=16
D17 VSS I DN AREA=2.037e-13 PJ=1.81e-06 $X=140 $Y=515 $D=32
.ENDS
***************************************
.SUBCKT ND3D3BWP7T A1 A2 A3 VDD ZN VSS
** N=8 EP=6 IP=0 FDC=18
M0 7 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 ZN A1 7 VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 7 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=2060 $Y=345 $D=0
M3 8 A2 7 VSS N L=1.8e-07 W=1e-06 $X=2780 $Y=345 $D=0
M4 7 A2 8 VSS N L=1.8e-07 W=1e-06 $X=3500 $Y=345 $D=0
M5 8 A2 7 VSS N L=1.8e-07 W=1e-06 $X=4220 $Y=345 $D=0
M6 VSS A3 8 VSS N L=1.8e-07 W=1e-06 $X=4940 $Y=345 $D=0
M7 8 A3 VSS VSS N L=1.8e-07 W=1e-06 $X=5660 $Y=345 $D=0
M8 VSS A3 8 VSS N L=1.8e-07 W=1e-06 $X=6380 $Y=345 $D=0
M9 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M10 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M11 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M12 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M13 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3500 $Y=2205 $D=16
M14 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4220 $Y=2205 $D=16
M15 ZN A3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4940 $Y=2205 $D=16
M16 VDD A3 ZN VDD P L=1.8e-07 W=1.37e-06 $X=5660 $Y=2205 $D=16
M17 ZN A3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=6380 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AN3D2BWP7T A1 A2 A3 Z VSS VDD
** N=9 EP=6 IP=0 FDC=10
M0 8 A1 7 VSS N L=1.8e-07 W=1e-06 $X=660 $Y=345 $D=0
M1 9 A2 8 VSS N L=1.8e-07 W=1e-06 $X=1380 $Y=345 $D=0
M2 VSS A3 9 VSS N L=1.8e-07 W=1e-06 $X=2100 $Y=345 $D=0
M3 Z 7 VSS VSS N L=1.8e-07 W=1e-06 $X=2820 $Y=345 $D=0
M4 VSS 7 Z VSS N L=1.8e-07 W=1e-06 $X=3540 $Y=345 $D=0
M5 VDD A1 7 VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M6 7 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1380 $Y=2205 $D=16
M7 VDD A3 7 VDD P L=1.8e-07 W=1.37e-06 $X=2100 $Y=2205 $D=16
M8 Z 7 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2820 $Y=2205 $D=16
M9 VDD 7 Z VDD P L=1.8e-07 W=1.37e-06 $X=3540 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OR3D2BWP7T A3 A2 A1 Z VDD VSS
** N=9 EP=6 IP=0 FDC=10
M0 VSS A3 7 VSS N L=1.8e-07 W=5e-07 $X=640 $Y=360 $D=0
M1 7 A2 VSS VSS N L=1.8e-07 W=5e-07 $X=1440 $Y=360 $D=0
M2 VSS A1 7 VSS N L=1.8e-07 W=5e-07 $X=2160 $Y=360 $D=0
M3 Z 7 VSS VSS N L=1.8e-07 W=1e-06 $X=2960 $Y=345 $D=0
M4 VSS 7 Z VSS N L=1.8e-07 W=1e-06 $X=3680 $Y=345 $D=0
M5 8 A3 7 VDD P L=1.8e-07 W=1.37e-06 $X=640 $Y=2205 $D=16
M6 9 A2 8 VDD P L=1.8e-07 W=1.37e-06 $X=1220 $Y=2205 $D=16
M7 VDD A1 9 VDD P L=1.8e-07 W=1.37e-06 $X=1800 $Y=2205 $D=16
M8 Z 7 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2600 $Y=2205 $D=16
M9 VDD 7 Z VDD P L=1.8e-07 W=1.37e-06 $X=3320 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT AOI32D1BWP7T A3 A2 A1 ZN B1 B2 VDD VSS
** N=12 EP=8 IP=0 FDC=10
M0 10 A3 VSS VSS N L=1.8e-07 W=1e-06 $X=680 $Y=345 $D=0
M1 11 A2 10 VSS N L=1.8e-07 W=1e-06 $X=1285 $Y=345 $D=0
M2 ZN A1 11 VSS N L=1.8e-07 W=1e-06 $X=1890 $Y=345 $D=0
M3 12 B1 ZN VSS N L=1.8e-07 W=1e-06 $X=2975 $Y=345 $D=0
M4 VSS B2 12 VSS N L=1.8e-07 W=1e-06 $X=3575 $Y=345 $D=0
M5 9 A3 ZN VDD P L=1.8e-07 W=1.37e-06 $X=680 $Y=2205 $D=16
M6 ZN A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=1400 $Y=2205 $D=16
M7 9 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2135 $Y=2205 $D=16
M8 VDD B1 9 VDD P L=1.8e-07 W=1.37e-06 $X=2855 $Y=2205 $D=16
M9 9 B2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3575 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ND4D3BWP7T A1 A2 A3 A4 VDD ZN VSS
** N=10 EP=7 IP=0 FDC=24
M0 8 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=665 $Y=345 $D=0
M1 ZN A1 8 VSS N L=1.8e-07 W=1e-06 $X=1385 $Y=345 $D=0
M2 8 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=2105 $Y=345 $D=0
M3 9 A2 8 VSS N L=1.8e-07 W=1e-06 $X=2825 $Y=345 $D=0
M4 8 A2 9 VSS N L=1.8e-07 W=1e-06 $X=3545 $Y=345 $D=0
M5 9 A2 8 VSS N L=1.8e-07 W=1e-06 $X=4265 $Y=345 $D=0
M6 10 A3 9 VSS N L=1.8e-07 W=1e-06 $X=4985 $Y=345 $D=0
M7 9 A3 10 VSS N L=1.8e-07 W=1e-06 $X=5705 $Y=345 $D=0
M8 10 A3 9 VSS N L=1.8e-07 W=1e-06 $X=6425 $Y=345 $D=0
M9 VSS A4 10 VSS N L=1.8e-07 W=1e-06 $X=7145 $Y=345 $D=0
M10 10 A4 VSS VSS N L=1.8e-07 W=1e-06 $X=7865 $Y=345 $D=0
M11 VSS A4 10 VSS N L=1.8e-07 W=1e-06 $X=8585 $Y=345 $D=0
M12 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=665 $Y=2205 $D=16
M13 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1385 $Y=2205 $D=16
M14 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2105 $Y=2205 $D=16
M15 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2825 $Y=2205 $D=16
M16 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3545 $Y=2205 $D=16
M17 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4265 $Y=2205 $D=16
M18 VDD A3 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4985 $Y=2205 $D=16
M19 ZN A3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=5705 $Y=2205 $D=16
M20 VDD A3 ZN VDD P L=1.8e-07 W=1.37e-06 $X=6425 $Y=2205 $D=16
M21 ZN A4 VDD VDD P L=1.8e-07 W=1.37e-06 $X=7145 $Y=2205 $D=16
M22 VDD A4 ZN VDD P L=1.8e-07 W=1.37e-06 $X=7865 $Y=2205 $D=16
M23 ZN A4 VDD VDD P L=1.8e-07 W=1.37e-06 $X=8585 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IND3D2BWP7T A1 VSS B1 B2 ZN VDD
** N=9 EP=6 IP=0 FDC=14
M0 VSS A1 7 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 8 7 VSS VSS N L=1.8e-07 W=1e-06 $X=1480 $Y=345 $D=0
M2 VSS 7 8 VSS N L=1.8e-07 W=1e-06 $X=2245 $Y=345 $D=0
M3 8 B1 9 VSS N L=1.8e-07 W=1e-06 $X=3665 $Y=345 $D=0
M4 9 B1 8 VSS N L=1.8e-07 W=1e-06 $X=4385 $Y=345 $D=0
M5 ZN B2 9 VSS N L=1.8e-07 W=1e-06 $X=5145 $Y=345 $D=0
M6 9 B2 ZN VSS N L=1.8e-07 W=1e-06 $X=5865 $Y=345 $D=0
M7 VDD A1 7 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M8 ZN 7 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1480 $Y=2205 $D=16
M9 VDD 7 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2245 $Y=2205 $D=16
M10 ZN B1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3665 $Y=2205 $D=16
M11 VDD B1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4385 $Y=2205 $D=16
M12 ZN B2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=5145 $Y=2205 $D=16
M13 VDD B2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=5865 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKND2D2BWP7T A2 VSS A1 ZN VDD
** N=6 EP=5 IP=0 FDC=8
M0 VSS A2 6 VSS N L=1.8e-07 W=6e-07 $X=660 $Y=545 $D=0
M1 6 A2 VSS VSS N L=1.8e-07 W=6e-07 $X=1380 $Y=545 $D=0
M2 ZN A1 6 VSS N L=1.8e-07 W=8e-07 $X=2320 $Y=545 $D=0
M3 6 A1 ZN VSS N L=1.8e-07 W=8e-07 $X=3120 $Y=545 $D=0
M4 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M5 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1380 $Y=2205 $D=16
M6 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2320 $Y=2205 $D=16
M7 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3120 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_24 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480
+ 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500
+ 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520
+ 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540
+ 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560
+ 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580
+ 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600
+ 601 602 603 604 605 606 607 608 609 610 611 612 613 614 616 617 618 619 620 621
+ 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729
** N=1395 EP=727 IP=6506 FDC=9928
M0 1381 989 230 1 N L=1.8e-07 W=9.05e-07 $X=107530 $Y=310425 $D=0
M1 1382 1032 1381 1 N L=1.8e-07 W=9.05e-07 $X=108130 $Y=310425 $D=0
M2 1 1039 1382 1 N L=1.8e-07 W=9.05e-07 $X=108730 $Y=310425 $D=0
M3 1383 1039 1 1 N L=1.8e-07 W=9.05e-07 $X=109600 $Y=310425 $D=0
M4 1384 1032 1383 1 N L=1.8e-07 W=9.05e-07 $X=110210 $Y=310425 $D=0
M5 230 989 1384 1 N L=1.8e-07 W=9.05e-07 $X=110820 $Y=310425 $D=0
M6 1385 1032 1 1 N L=1.8e-07 W=1e-06 $X=112470 $Y=310425 $D=0
M7 230 992 1385 1 N L=1.8e-07 W=1e-06 $X=113070 $Y=310425 $D=0
M8 1386 992 230 1 N L=1.8e-07 W=1e-06 $X=113790 $Y=310425 $D=0
M9 1 1032 1386 1 N L=1.8e-07 W=1e-06 $X=114395 $Y=310425 $D=0
M10 1387 1082 1092 1 N L=1.8e-07 W=1e-06 $X=135440 $Y=310425 $D=0
M11 1388 1085 1387 1 N L=1.8e-07 W=1e-06 $X=136160 $Y=310425 $D=0
M12 1389 260 1388 1 N L=1.8e-07 W=1e-06 $X=136880 $Y=310425 $D=0
M13 1 957 1389 1 N L=1.8e-07 W=1e-06 $X=137600 $Y=310425 $D=0
M14 265 1092 1 1 N L=1.8e-07 W=1e-06 $X=138320 $Y=310425 $D=0
M15 1 1092 265 1 N L=1.8e-07 W=1e-06 $X=139040 $Y=310425 $D=0
M16 1390 1047 1 1 N L=1.8e-07 W=5e-07 $X=146665 $Y=308970 $D=0
M17 1391 1072 1390 1 N L=1.8e-07 W=5e-07 $X=147275 $Y=308970 $D=0
M18 1105 281 1391 1 N L=1.8e-07 W=5e-07 $X=147885 $Y=308970 $D=0
M19 1392 280 1105 1 N L=1.8e-07 W=5e-07 $X=148965 $Y=308970 $D=0
M20 1 1072 1392 1 N L=1.8e-07 W=5e-07 $X=149565 $Y=308970 $D=0
M21 1158 340 1 1 N L=1.8e-07 W=8e-07 $X=207865 $Y=324520 $D=0
M22 1160 1158 1 1 N L=1.8e-07 W=8.3e-07 $X=209385 $Y=324490 $D=0
M23 1 1158 1160 1 N L=1.8e-07 W=8.3e-07 $X=210105 $Y=324490 $D=0
M24 1393 1355 1 1 N L=1.8e-07 W=1e-06 $X=446240 $Y=294745 $D=0
M25 1167 661 1393 1 N L=1.8e-07 W=1e-06 $X=446960 $Y=294745 $D=0
M26 1394 661 1167 1 N L=1.8e-07 W=1e-06 $X=447680 $Y=294745 $D=0
M27 1 1355 1394 1 N L=1.8e-07 W=1e-06 $X=448400 $Y=294745 $D=0
M28 1395 524 1 1 N L=1.8e-07 W=1e-06 $X=449240 $Y=294745 $D=0
M29 1355 1359 1395 1 N L=1.8e-07 W=1e-06 $X=449840 $Y=294745 $D=0
M30 230 1032 1052 2 P L=1.8e-07 W=1.275e-06 $X=107490 $Y=312380 $D=16
M31 1052 1032 230 2 P L=1.8e-07 W=1.275e-06 $X=108210 $Y=312380 $D=16
M32 230 1039 1052 2 P L=1.8e-07 W=1.275e-06 $X=109030 $Y=312380 $D=16
M33 1052 1039 230 2 P L=1.8e-07 W=1.275e-06 $X=109750 $Y=312380 $D=16
M34 230 989 1052 2 P L=1.8e-07 W=1.275e-06 $X=110550 $Y=312380 $D=16
M35 1052 989 230 2 P L=1.8e-07 W=1.275e-06 $X=111270 $Y=312380 $D=16
M36 2 1032 1052 2 P L=1.8e-07 W=1.37e-06 $X=112230 $Y=312285 $D=16
M37 1052 992 2 2 P L=1.8e-07 W=1.37e-06 $X=112950 $Y=312285 $D=16
M38 2 992 1052 2 P L=1.8e-07 W=1.37e-06 $X=113670 $Y=312285 $D=16
M39 1052 1032 2 2 P L=1.8e-07 W=1.37e-06 $X=114395 $Y=312285 $D=16
M40 1092 1082 2 2 P L=1.8e-07 W=1.37e-06 $X=135440 $Y=312285 $D=16
M41 2 1085 1092 2 P L=1.8e-07 W=1.37e-06 $X=136160 $Y=312285 $D=16
M42 1092 260 2 2 P L=1.8e-07 W=1.37e-06 $X=136880 $Y=312285 $D=16
M43 2 957 1092 2 P L=1.8e-07 W=1.37e-06 $X=137600 $Y=312285 $D=16
M44 265 1092 2 2 P L=1.8e-07 W=1.37e-06 $X=138320 $Y=312285 $D=16
M45 2 1092 265 2 P L=1.8e-07 W=1.37e-06 $X=139040 $Y=312285 $D=16
M46 1107 1047 1105 2 P L=1.8e-07 W=6.85e-07 $X=146665 $Y=306915 $D=16
M47 1105 1072 1107 2 P L=1.8e-07 W=6.85e-07 $X=147390 $Y=306915 $D=16
M48 1107 281 1105 2 P L=1.8e-07 W=6.85e-07 $X=148125 $Y=306915 $D=16
M49 2 280 1107 2 P L=1.8e-07 W=6.85e-07 $X=148845 $Y=306915 $D=16
M50 1107 1072 2 2 P L=1.8e-07 W=6.85e-07 $X=149680 $Y=306915 $D=16
M51 1158 340 2 2 P L=1.8e-07 W=1.14e-06 $X=207140 $Y=322185 $D=16
M52 2 340 1158 2 P L=1.8e-07 W=1.14e-06 $X=207865 $Y=322185 $D=16
M53 1160 1158 2 2 P L=1.8e-07 W=1.37e-06 $X=208585 $Y=322185 $D=16
M54 2 1158 1160 2 P L=1.8e-07 W=1.37e-06 $X=209305 $Y=322185 $D=16
M55 1160 1158 2 2 P L=1.8e-07 W=1.37e-06 $X=210105 $Y=322185 $D=16
M56 1167 1355 2 2 P L=1.8e-07 W=1.37e-06 $X=446240 $Y=296605 $D=16
M57 2 661 1167 2 P L=1.8e-07 W=1.37e-06 $X=446960 $Y=296605 $D=16
M58 1167 661 2 2 P L=1.8e-07 W=1.37e-06 $X=447680 $Y=296605 $D=16
M59 2 1355 1167 2 P L=1.8e-07 W=1.37e-06 $X=448400 $Y=296605 $D=16
M60 1355 524 2 2 P L=1.8e-07 W=1.37e-06 $X=449120 $Y=296605 $D=16
M61 2 1359 1355 2 P L=1.8e-07 W=1.37e-06 $X=449840 $Y=296605 $D=16
D62 1 340 DN AREA=2.037e-13 PJ=1.81e-06 $X=206620 $Y=324420 $D=32
X148 1 605 ANTENNABWP7T $T=474160 302240 0 180 $X=472750 $Y=298030
X149 1 675 ANTENNABWP7T $T=474160 310080 0 180 $X=472750 $Y=305870
X150 1 678 ANTENNABWP7T $T=473040 310080 0 0 $X=472750 $Y=309845
X151 1 600 ANTENNABWP7T $T=474160 317920 0 180 $X=472750 $Y=313710
X152 1 707 ANTENNABWP7T $T=473040 317920 0 0 $X=472750 $Y=317685
X153 1 690 ANTENNABWP7T $T=474160 325760 0 180 $X=472750 $Y=321550
X154 1 724 ANTENNABWP7T $T=473040 325760 0 0 $X=472750 $Y=325525
X155 1 727 ANTENNABWP7T $T=474160 333600 0 180 $X=472750 $Y=329390
X156 1 449 ANTENNABWP7T $T=473040 333600 0 0 $X=472750 $Y=333365
X157 1 684 ANTENNABWP7T $T=474160 341440 0 180 $X=472750 $Y=337230
X158 1 728 ANTENNABWP7T $T=474160 349280 0 180 $X=472750 $Y=345070
X159 1 630 ANTENNABWP7T $T=473040 349280 0 0 $X=472750 $Y=349045
X160 1 697 ANTENNABWP7T $T=474160 357120 0 180 $X=472750 $Y=352910
X161 1 701 712 ICV_1 $T=469680 294400 0 0 $X=469390 $Y=294165
X162 1 492 617 ICV_1 $T=469680 302240 0 0 $X=469390 $Y=302005
X163 1 500 529 ICV_1 $T=469680 341440 0 0 $X=469390 $Y=341205
X164 1 518 686 ICV_1 $T=470800 310080 0 0 $X=470510 $Y=309845
X165 1 635 514 ICV_1 $T=470800 317920 0 0 $X=470510 $Y=317685
X166 1 715 716 ICV_1 $T=470800 325760 0 0 $X=470510 $Y=325525
X167 1 708 677 ICV_1 $T=470800 333600 0 0 $X=470510 $Y=333365
X168 1 709 718 ICV_1 $T=470800 349280 0 0 $X=470510 $Y=349045
X169 1 637 725 ICV_1 $T=471920 294400 0 0 $X=471630 $Y=294165
X170 1 729 726 ICV_1 $T=471920 302240 0 0 $X=471630 $Y=302005
X171 1 717 458 ICV_1 $T=471920 341440 0 0 $X=471630 $Y=341205
X172 1 720 713 ICV_2 $T=471920 302240 0 180 $X=470510 $Y=298030
X173 1 591 485 ICV_2 $T=471920 310080 0 180 $X=470510 $Y=305870
X174 1 705 710 ICV_2 $T=471920 317920 0 180 $X=470510 $Y=313710
X175 1 721 714 ICV_2 $T=471920 325760 0 180 $X=470510 $Y=321550
X176 1 722 711 ICV_2 $T=471920 333600 0 180 $X=470510 $Y=329390
X177 1 719 490 ICV_2 $T=471920 341440 0 180 $X=470510 $Y=337230
X178 1 585 440 ICV_2 $T=471920 349280 0 180 $X=470510 $Y=345070
X179 1 723 670 ICV_2 $T=471920 357120 0 180 $X=470510 $Y=352910
X262 19 1 2 869 CKBD1BWP7T $T=24480 325760 0 0 $X=24190 $Y=325525
X263 1053 1 2 277 CKBD1BWP7T $T=139840 317920 1 0 $X=139550 $Y=313710
X264 1090 1 2 282 CKBD1BWP7T $T=146000 294400 0 0 $X=145710 $Y=294165
X265 1104 1 2 288 CKBD1BWP7T $T=151600 310080 0 0 $X=151310 $Y=309845
X266 1051 1 2 291 CKBD1BWP7T $T=153840 310080 0 0 $X=153550 $Y=309845
X267 1087 1 2 1112 CKBD1BWP7T $T=154400 317920 0 0 $X=154110 $Y=317685
X268 1097 1 2 293 CKBD1BWP7T $T=154400 325760 1 0 $X=154110 $Y=321550
X269 300 1 2 302 CKBD1BWP7T $T=168400 357120 1 0 $X=168110 $Y=352910
X270 306 1 2 309 CKBD1BWP7T $T=174000 357120 1 0 $X=173710 $Y=352910
X271 341 1 2 344 CKBD1BWP7T $T=206480 310080 0 0 $X=206190 $Y=309845
X272 343 1 2 347 CKBD1BWP7T $T=207040 349280 1 0 $X=206750 $Y=345070
X273 1168 1 2 360 CKBD1BWP7T $T=218800 325760 1 0 $X=218510 $Y=321550
X274 1170 1 2 364 CKBD1BWP7T $T=219920 302240 0 0 $X=219630 $Y=302005
X275 1172 1 2 374 CKBD1BWP7T $T=236720 341440 0 180 $X=234190 $Y=337230
X276 1182 1 2 373 CKBD1BWP7T $T=237840 349280 1 180 $X=235310 $Y=349045
X277 1178 1 2 386 CKBD1BWP7T $T=238400 341440 1 0 $X=238110 $Y=337230
X278 1208 1 2 413 CKBD1BWP7T $T=263040 310080 1 0 $X=262750 $Y=305870
X279 417 1 2 1173 CKBD1BWP7T $T=269200 310080 0 180 $X=266670 $Y=305870
X280 1217 1 2 1136 CKBD1BWP7T $T=273120 333600 0 180 $X=270590 $Y=329390
X281 471 1 2 1216 CKBD1BWP7T $T=310080 325760 0 180 $X=307550 $Y=321550
X282 490 1 2 488 CKBD1BWP7T $T=316240 317920 0 180 $X=313710 $Y=313710
X283 492 1 2 457 CKBD1BWP7T $T=318480 302240 0 180 $X=315950 $Y=298030
X284 529 1 2 527 CKBD1BWP7T $T=346480 341440 1 180 $X=343950 $Y=341205
X285 532 1 2 1282 CKBD1BWP7T $T=347040 333600 1 0 $X=346750 $Y=329390
X286 534 1 2 533 CKBD1BWP7T $T=349280 341440 0 180 $X=346750 $Y=337230
X287 1299 1 2 543 CKBD1BWP7T $T=364960 302240 0 180 $X=362430 $Y=298030
X288 565 1 2 564 CKBD1BWP7T $T=378960 325760 0 180 $X=376430 $Y=321550
X289 565 1 2 567 CKBD1BWP7T $T=381200 325760 0 180 $X=378670 $Y=321550
X290 585 1 2 583 CKBD1BWP7T $T=389600 317920 1 180 $X=387070 $Y=317685
X291 600 1 2 515 CKBD1BWP7T $T=400800 325760 1 180 $X=398270 $Y=325525
X292 580 1 2 562 CKBD1BWP7T $T=408080 325760 1 180 $X=405550 $Y=325525
X293 1338 1 2 616 CKBD1BWP7T $T=421520 302240 1 180 $X=418990 $Y=302005
X294 376 1 2 658 CKBD1BWP7T $T=443920 333600 1 0 $X=443630 $Y=329390
X295 617 1 2 674 CKBD1BWP7T $T=460160 325760 0 0 $X=459870 $Y=325525
X296 635 1 2 698 CKBD1BWP7T $T=470800 349280 0 180 $X=468270 $Y=345070
X297 873 1 2 887 INVD0BWP7T $T=39040 341440 0 0 $X=38750 $Y=341205
X298 45 1 2 890 INVD0BWP7T $T=39600 310080 1 0 $X=39310 $Y=305870
X299 54 1 2 875 INVD0BWP7T $T=43520 310080 1 180 $X=41550 $Y=309845
X300 896 1 2 913 INVD0BWP7T $T=48000 325760 1 0 $X=47710 $Y=321550
X301 81 1 2 906 INVD0BWP7T $T=50240 341440 1 180 $X=48270 $Y=341205
X302 928 1 2 925 INVD0BWP7T $T=55840 310080 1 0 $X=55550 $Y=305870
X303 9 1 2 935 INVD0BWP7T $T=58640 310080 0 0 $X=58350 $Y=309845
X304 46 1 2 983 INVD0BWP7T $T=79920 341440 1 0 $X=79630 $Y=337230
X305 171 1 2 969 INVD0BWP7T $T=87760 349280 1 180 $X=85790 $Y=349045
X306 989 1 2 159 INVD0BWP7T $T=88880 310080 0 180 $X=86910 $Y=305870
X307 991 1 2 977 INVD0BWP7T $T=91680 333600 0 180 $X=89710 $Y=329390
X308 990 1 2 187 INVD0BWP7T $T=91680 310080 1 0 $X=91390 $Y=305870
X309 100 1 2 190 INVD0BWP7T $T=95040 317920 0 180 $X=93070 $Y=313710
X310 229 1 2 1020 INVD0BWP7T $T=112960 302240 0 180 $X=110990 $Y=298030
X311 913 1 2 1056 INVD0BWP7T $T=121920 317920 1 0 $X=121630 $Y=313710
X312 1045 1 2 1004 INVD0BWP7T $T=128080 325760 0 180 $X=126110 $Y=321550
X313 252 1 2 1025 INVD0BWP7T $T=132000 333600 1 180 $X=130030 $Y=333365
X314 1054 1 2 1084 INVD0BWP7T $T=133120 325760 1 0 $X=132830 $Y=321550
X315 1083 1 2 1086 INVD0BWP7T $T=134800 325760 0 0 $X=134510 $Y=325525
X316 1089 1 2 1074 INVD0BWP7T $T=136480 341440 1 180 $X=134510 $Y=341205
X317 945 1 2 1094 INVD0BWP7T $T=137600 317920 0 0 $X=137310 $Y=317685
X318 914 1 2 1096 INVD0BWP7T $T=138160 333600 1 0 $X=137870 $Y=329390
X319 911 1 2 1078 INVD0BWP7T $T=138720 325760 0 0 $X=138430 $Y=325525
X320 927 1 2 280 INVD0BWP7T $T=144320 302240 0 0 $X=144030 $Y=302005
X321 1109 1 2 1100 INVD0BWP7T $T=150480 341440 0 180 $X=148510 $Y=337230
X322 1111 1 2 1013 INVD0BWP7T $T=152720 341440 0 180 $X=150750 $Y=337230
X323 294 1 2 1113 INVD0BWP7T $T=163920 302240 1 0 $X=163630 $Y=298030
X324 277 1 2 297 INVD0BWP7T $T=163920 310080 1 0 $X=163630 $Y=305870
X325 293 1 2 1117 INVD0BWP7T $T=165600 310080 1 0 $X=165310 $Y=305870
X326 1112 1 2 1114 INVD0BWP7T $T=167840 317920 0 0 $X=167550 $Y=317685
X327 285 1 2 1122 INVD0BWP7T $T=169520 349280 0 0 $X=169230 $Y=349045
X328 1115 1 2 1129 INVD0BWP7T $T=173440 333600 1 0 $X=173150 $Y=329390
X329 378 1 2 380 INVD0BWP7T $T=233920 317920 1 0 $X=233630 $Y=313710
X330 442 1 2 1232 INVD0BWP7T $T=281520 302240 1 0 $X=281230 $Y=298030
X331 1186 1 2 1241 INVD0BWP7T $T=293280 325760 1 0 $X=292990 $Y=321550
X332 471 1 2 1218 INVD0BWP7T $T=304480 325760 0 180 $X=302510 $Y=321550
X333 1253 1 2 1240 INVD0BWP7T $T=304480 341440 0 180 $X=302510 $Y=337230
X334 519 1 2 1275 INVD0BWP7T $T=340320 317920 1 180 $X=338350 $Y=317685
X335 1278 1 2 1286 INVD0BWP7T $T=345360 333600 0 0 $X=345070 $Y=333365
X336 532 1 2 1281 INVD0BWP7T $T=348160 325760 1 180 $X=346190 $Y=325525
X337 1291 1 2 1284 INVD0BWP7T $T=354320 302240 0 180 $X=352350 $Y=298030
X338 1298 1 2 1305 INVD0BWP7T $T=364400 325760 0 0 $X=364110 $Y=325525
X339 580 1 2 1313 INVD0BWP7T $T=386240 341440 0 180 $X=384270 $Y=337230
X340 1323 1 2 1320 INVD0BWP7T $T=391840 333600 0 180 $X=389870 $Y=329390
X341 1331 1 2 1333 INVD0BWP7T $T=417040 333600 0 0 $X=416750 $Y=333365
X342 1336 1 2 627 INVD0BWP7T $T=424320 357120 1 0 $X=424030 $Y=352910
X343 649 1 2 1353 INVD0BWP7T $T=450640 325760 0 180 $X=448670 $Y=321550
X344 1148 1 2 1356 INVD0BWP7T $T=449520 317920 1 0 $X=449230 $Y=313710
X345 384 1 2 1358 INVD0BWP7T $T=457920 341440 0 0 $X=457630 $Y=341205
X346 1354 1 2 1364 INVD0BWP7T $T=461280 341440 0 0 $X=460990 $Y=341205
X347 326 1 2 1361 INVD0BWP7T $T=463520 310080 1 0 $X=463230 $Y=305870
X348 684 1 2 1357 INVD0BWP7T $T=465200 333600 1 180 $X=463230 $Y=333365
X349 487 1 2 1362 INVD0BWP7T $T=467440 294400 1 180 $X=465470 $Y=294165
X350 1095 286 1 2 BUFFD1P5BWP7T $T=148800 294400 0 0 $X=148510 $Y=294165
X351 1140 349 1 2 BUFFD1P5BWP7T $T=207040 310080 1 0 $X=206750 $Y=305870
X352 354 355 1 2 BUFFD1P5BWP7T $T=213760 357120 1 0 $X=213470 $Y=352910
X353 1128 359 1 2 BUFFD1P5BWP7T $T=216000 317920 0 0 $X=215710 $Y=317685
X354 485 483 1 2 BUFFD1P5BWP7T $T=312880 302240 1 180 $X=309790 $Y=302005
X355 493 1133 1 2 BUFFD1P5BWP7T $T=318480 357120 0 180 $X=315390 $Y=352910
X356 503 468 1 2 BUFFD1P5BWP7T $T=324640 357120 0 180 $X=321550 $Y=352910
X357 514 511 1 2 BUFFD1P5BWP7T $T=338640 325760 0 180 $X=335550 $Y=321550
X358 1318 569 1 2 BUFFD1P5BWP7T $T=382320 310080 0 180 $X=379230 $Y=305870
X359 591 590 1 2 BUFFD1P5BWP7T $T=395200 310080 0 180 $X=392110 $Y=305870
X360 605 601 1 2 BUFFD1P5BWP7T $T=404720 302240 0 180 $X=401630 $Y=298030
X361 637 432 1 2 BUFFD1P5BWP7T $T=437760 333600 0 180 $X=434670 $Y=329390
X362 1350 509 1 2 BUFFD1P5BWP7T $T=440000 317920 0 180 $X=436910 $Y=313710
X363 678 673 1 2 BUFFD1P5BWP7T $T=465200 317920 0 180 $X=462110 $Y=313710
X364 691 462 1 2 BUFFD1P5BWP7T $T=468560 349280 0 180 $X=465470 $Y=345070
X365 697 682 1 2 BUFFD1P5BWP7T $T=469680 341440 1 180 $X=466590 $Y=341205
X366 700 693 1 2 BUFFD1P5BWP7T $T=470240 333600 1 180 $X=467150 $Y=333365
X367 702 425 1 2 BUFFD1P5BWP7T $T=470800 302240 0 180 $X=467710 $Y=298030
X368 703 443 1 2 BUFFD1P5BWP7T $T=470800 341440 0 180 $X=467710 $Y=337230
X369 704 694 1 2 BUFFD1P5BWP7T $T=470800 357120 0 180 $X=467710 $Y=352910
X370 410 1202 2 1 397 1212 1206 MAOI22D0BWP7T $T=261360 333600 0 0 $X=261070 $Y=333365
X371 421 422 2 1 397 1214 1221 MAOI22D0BWP7T $T=270320 341440 1 0 $X=270030 $Y=337230
X372 444 449 2 1 449 1224 444 MAOI22D0BWP7T $T=283200 333600 0 180 $X=278990 $Y=329390
X373 581 670 2 1 581 1359 670 MAOI22D0BWP7T $T=465200 302240 0 180 $X=460990 $Y=298030
X448 272 1115 299 272 1 1115 2 IAO22D2BWP7T $T=163920 333600 1 0 $X=163630 $Y=329390
X449 324 286 1146 324 1 286 2 IAO22D2BWP7T $T=197520 302240 1 180 $X=191070 $Y=302005
X450 458 1218 1243 458 1 1218 2 IAO22D2BWP7T $T=293280 333600 0 0 $X=292990 $Y=333365
X451 577 1313 1315 577 1 1313 2 IAO22D2BWP7T $T=389600 357120 0 180 $X=383150 $Y=352910
X452 895 1 2 892 BUFFD1BWP7T $T=43520 325760 0 180 $X=40990 $Y=321550
X453 882 1 2 902 BUFFD1BWP7T $T=43520 325760 1 0 $X=43230 $Y=321550
X454 923 1 2 957 BUFFD1BWP7T $T=62000 325760 1 0 $X=61710 $Y=321550
X455 1001 1 2 1011 BUFFD1BWP7T $T=93360 333600 0 0 $X=93070 $Y=333365
X456 1012 1 2 1010 BUFFD1BWP7T $T=97840 310080 0 180 $X=95310 $Y=305870
X457 162 1 2 1017 BUFFD1BWP7T $T=98960 341440 0 0 $X=98670 $Y=341205
X458 1026 1 2 1021 BUFFD1BWP7T $T=102880 310080 1 180 $X=100350 $Y=309845
X459 1014 1 2 1035 BUFFD1BWP7T $T=102880 333600 0 0 $X=102590 $Y=333365
X460 933 1 2 1058 BUFFD1BWP7T $T=121920 325760 0 0 $X=121630 $Y=325525
X461 929 1 2 238 BUFFD1BWP7T $T=122480 310080 0 0 $X=122190 $Y=309845
X462 988 1 2 1064 BUFFD1BWP7T $T=124720 317920 1 0 $X=124430 $Y=313710
X463 1003 1 2 1073 BUFFD1BWP7T $T=128080 333600 0 0 $X=127790 $Y=333365
X464 253 1 2 1080 BUFFD1BWP7T $T=130880 349280 0 0 $X=130590 $Y=349045
X465 1081 1 2 1088 BUFFD1BWP7T $T=134240 341440 1 0 $X=133950 $Y=337230
X466 1068 1 2 1091 BUFFD1BWP7T $T=135920 333600 1 0 $X=135630 $Y=329390
X467 1008 1 2 1103 BUFFD1BWP7T $T=144320 325760 1 0 $X=144030 $Y=321550
X468 1105 1 2 284 BUFFD1BWP7T $T=148240 302240 0 0 $X=147950 $Y=302005
X469 1075 1 2 1115 BUFFD1BWP7T $T=170080 333600 1 0 $X=169790 $Y=329390
X470 358 1 2 1163 BUFFD1BWP7T $T=217680 294400 0 0 $X=217390 $Y=294165
X471 475 1 2 477 BUFFD1BWP7T $T=305600 357120 1 0 $X=305310 $Y=352910
X472 519 1 2 505 BUFFD1BWP7T $T=340320 317920 0 0 $X=340030 $Y=317685
X473 1283 1 2 1217 BUFFD1BWP7T $T=343120 333600 0 180 $X=340590 $Y=329390
X474 537 1 2 536 BUFFD1BWP7T $T=353760 294400 1 180 $X=351230 $Y=294165
X475 1307 1 2 1169 BUFFD1BWP7T $T=367200 310080 0 180 $X=364670 $Y=305870
X476 1308 1 2 1302 BUFFD1BWP7T $T=367200 333600 1 180 $X=364670 $Y=333365
X477 331 1 2 570 BUFFD1BWP7T $T=377840 325760 0 0 $X=377550 $Y=325525
X478 609 1 2 608 BUFFD1BWP7T $T=406960 310080 1 180 $X=404430 $Y=309845
X479 1335 1 2 618 BUFFD1BWP7T $T=418720 341440 1 0 $X=418430 $Y=337230
X480 619 1 2 1337 BUFFD1BWP7T $T=419840 302240 1 0 $X=419550 $Y=298030
X481 648 1 2 643 BUFFD1BWP7T $T=443920 333600 1 180 $X=441390 $Y=333365
X482 375 1 2 663 BUFFD1BWP7T $T=448960 341440 0 0 $X=448670 $Y=341205
X483 1360 1 2 671 BUFFD1BWP7T $T=460720 349280 0 0 $X=460430 $Y=349045
X484 602 1 2 1354 BUFFD1BWP7T $T=463520 310080 0 180 $X=460990 $Y=305870
X485 1363 1 2 680 BUFFD1BWP7T $T=462960 333600 1 0 $X=462670 $Y=329390
X486 1 2 DCAP4BWP7T $T=39600 349280 1 0 $X=39310 $Y=345070
X487 1 2 DCAP4BWP7T $T=45760 325760 1 0 $X=45470 $Y=321550
X488 1 2 DCAP4BWP7T $T=124160 325760 0 0 $X=123870 $Y=325525
X489 1 2 DCAP4BWP7T $T=124720 310080 0 0 $X=124430 $Y=309845
X490 1 2 DCAP4BWP7T $T=136480 325760 0 0 $X=136190 $Y=325525
X491 1 2 DCAP4BWP7T $T=138720 302240 0 0 $X=138430 $Y=302005
X492 1 2 DCAP4BWP7T $T=139840 310080 1 0 $X=139550 $Y=305870
X493 1 2 DCAP4BWP7T $T=139840 310080 0 0 $X=139550 $Y=309845
X494 1 2 DCAP4BWP7T $T=152160 317920 0 0 $X=151870 $Y=317685
X495 1 2 DCAP4BWP7T $T=209840 310080 1 0 $X=209550 $Y=305870
X496 1 2 DCAP4BWP7T $T=213760 349280 1 0 $X=213470 $Y=345070
X497 1 2 DCAP4BWP7T $T=273680 317920 0 0 $X=273390 $Y=317685
X498 1 2 DCAP4BWP7T $T=283760 317920 1 0 $X=283470 $Y=313710
X499 1 2 DCAP4BWP7T $T=296080 349280 0 0 $X=295790 $Y=349045
X500 1 2 DCAP4BWP7T $T=296080 357120 1 0 $X=295790 $Y=352910
X501 1 2 DCAP4BWP7T $T=303920 310080 0 0 $X=303630 $Y=309845
X502 1 2 DCAP4BWP7T $T=342560 317920 0 0 $X=342270 $Y=317685
X503 1 2 DCAP4BWP7T $T=348720 317920 1 0 $X=348430 $Y=313710
X504 1 2 DCAP4BWP7T $T=377840 333600 1 0 $X=377550 $Y=329390
X505 1 2 DCAP4BWP7T $T=380080 341440 0 0 $X=379790 $Y=341205
X506 1 2 DCAP4BWP7T $T=395200 341440 0 0 $X=394910 $Y=341205
X507 1 2 DCAP4BWP7T $T=422080 357120 1 0 $X=421790 $Y=352910
X508 1 2 DCAP4BWP7T $T=431040 333600 1 0 $X=430750 $Y=329390
X509 1 2 DCAP4BWP7T $T=433840 325760 0 0 $X=433550 $Y=325525
X510 1 2 DCAP4BWP7T $T=465200 310080 1 0 $X=464910 $Y=305870
X511 1 2 DCAP4BWP7T $T=465760 341440 1 0 $X=465470 $Y=337230
X512 1 2 ICV_3 $T=31200 302240 0 0 $X=30910 $Y=302005
X513 1 2 ICV_3 $T=31200 325760 0 0 $X=30910 $Y=325525
X514 1 2 ICV_3 $T=31200 333600 1 0 $X=30910 $Y=329390
X515 1 2 ICV_3 $T=31200 333600 0 0 $X=30910 $Y=333365
X516 1 2 ICV_3 $T=31200 349280 1 0 $X=30910 $Y=345070
X517 1 2 ICV_3 $T=31200 349280 0 0 $X=30910 $Y=349045
X518 1 2 ICV_3 $T=73200 333600 1 0 $X=72910 $Y=329390
X519 1 2 ICV_3 $T=96720 349280 1 0 $X=96430 $Y=345070
X520 1 2 ICV_3 $T=98400 302240 1 0 $X=98110 $Y=298030
X521 1 2 ICV_3 $T=98400 341440 1 0 $X=98110 $Y=337230
X522 1 2 ICV_3 $T=115200 310080 0 0 $X=114910 $Y=309845
X523 1 2 ICV_3 $T=119120 325760 0 0 $X=118830 $Y=325525
X524 1 2 ICV_3 $T=133120 349280 0 0 $X=132830 $Y=349045
X525 1 2 ICV_3 $T=143200 294400 0 0 $X=142910 $Y=294165
X526 1 2 ICV_3 $T=157200 294400 0 0 $X=156910 $Y=294165
X527 1 2 ICV_3 $T=157200 302240 0 0 $X=156910 $Y=302005
X528 1 2 ICV_3 $T=157200 325760 0 0 $X=156910 $Y=325525
X529 1 2 ICV_3 $T=157200 333600 0 0 $X=156910 $Y=333365
X530 1 2 ICV_3 $T=181280 317920 1 0 $X=180990 $Y=313710
X531 1 2 ICV_3 $T=181280 333600 0 0 $X=180990 $Y=333365
X532 1 2 ICV_3 $T=182960 325760 1 0 $X=182670 $Y=321550
X533 1 2 ICV_3 $T=199200 294400 0 0 $X=198910 $Y=294165
X534 1 2 ICV_3 $T=199200 310080 1 0 $X=198910 $Y=305870
X535 1 2 ICV_3 $T=199200 325760 1 0 $X=198910 $Y=321550
X536 1 2 ICV_3 $T=199200 325760 0 0 $X=198910 $Y=325525
X537 1 2 ICV_3 $T=226640 317920 0 0 $X=226350 $Y=317685
X538 1 2 ICV_3 $T=241200 357120 1 0 $X=240910 $Y=352910
X539 1 2 ICV_3 $T=249600 310080 1 0 $X=249310 $Y=305870
X540 1 2 ICV_3 $T=269200 310080 1 0 $X=268910 $Y=305870
X541 1 2 ICV_3 $T=287120 333600 1 0 $X=286830 $Y=329390
X542 1 2 ICV_3 $T=291600 341440 0 0 $X=291310 $Y=341205
X543 1 2 ICV_3 $T=302800 357120 1 0 $X=302510 $Y=352910
X544 1 2 ICV_3 $T=325200 294400 0 0 $X=324910 $Y=294165
X545 1 2 ICV_3 $T=325200 317920 1 0 $X=324910 $Y=313710
X546 1 2 ICV_3 $T=333600 317920 1 0 $X=333310 $Y=313710
X547 1 2 ICV_3 $T=338080 333600 1 0 $X=337790 $Y=329390
X548 1 2 ICV_3 $T=367200 310080 1 0 $X=366910 $Y=305870
X549 1 2 ICV_3 $T=367200 310080 0 0 $X=366910 $Y=309845
X550 1 2 ICV_3 $T=367200 333600 0 0 $X=366910 $Y=333365
X551 1 2 ICV_3 $T=367200 357120 1 0 $X=366910 $Y=352910
X552 1 2 ICV_3 $T=375600 317920 1 0 $X=375310 $Y=313710
X553 1 2 ICV_3 $T=380080 325760 0 0 $X=379790 $Y=325525
X554 1 2 ICV_3 $T=409200 317920 0 0 $X=408910 $Y=317685
X555 1 2 ICV_3 $T=436080 310080 1 0 $X=435790 $Y=305870
X556 1 2 ICV_3 $T=442800 294400 0 0 $X=442510 $Y=294165
X557 1 2 ICV_3 $T=451200 341440 0 0 $X=450910 $Y=341205
X558 1 2 DCAP8BWP7T $T=26160 310080 0 0 $X=25870 $Y=309845
X559 1 2 DCAP8BWP7T $T=28960 302240 1 0 $X=28670 $Y=298030
X560 1 2 DCAP8BWP7T $T=29520 357120 1 0 $X=29230 $Y=352910
X561 1 2 DCAP8BWP7T $T=35120 317920 1 0 $X=34830 $Y=313710
X562 1 2 DCAP8BWP7T $T=44080 349280 0 0 $X=43790 $Y=349045
X563 1 2 DCAP8BWP7T $T=112960 294400 0 0 $X=112670 $Y=294165
X564 1 2 DCAP8BWP7T $T=129200 341440 1 0 $X=128910 $Y=337230
X565 1 2 DCAP8BWP7T $T=139280 349280 0 0 $X=138990 $Y=349045
X566 1 2 DCAP8BWP7T $T=146560 325760 1 0 $X=146270 $Y=321550
X567 1 2 DCAP8BWP7T $T=150480 310080 1 0 $X=150190 $Y=305870
X568 1 2 DCAP8BWP7T $T=155520 333600 1 0 $X=155230 $Y=329390
X569 1 2 DCAP8BWP7T $T=155520 349280 0 0 $X=155230 $Y=349045
X570 1 2 DCAP8BWP7T $T=165600 325760 1 0 $X=165310 $Y=321550
X571 1 2 DCAP8BWP7T $T=171200 349280 0 0 $X=170910 $Y=349045
X572 1 2 DCAP8BWP7T $T=176240 357120 1 0 $X=175950 $Y=352910
X573 1 2 DCAP8BWP7T $T=188000 349280 0 0 $X=187710 $Y=349045
X574 1 2 DCAP8BWP7T $T=196960 341440 1 0 $X=196670 $Y=337230
X575 1 2 DCAP8BWP7T $T=197520 302240 0 0 $X=197230 $Y=302005
X576 1 2 DCAP8BWP7T $T=197520 317920 1 0 $X=197230 $Y=313710
X577 1 2 DCAP8BWP7T $T=216560 357120 1 0 $X=216270 $Y=352910
X578 1 2 DCAP8BWP7T $T=217120 325760 0 0 $X=216830 $Y=325525
X579 1 2 DCAP8BWP7T $T=221600 317920 1 0 $X=221310 $Y=313710
X580 1 2 DCAP8BWP7T $T=236160 325760 1 0 $X=235870 $Y=321550
X581 1 2 DCAP8BWP7T $T=239520 333600 0 0 $X=239230 $Y=333365
X582 1 2 DCAP8BWP7T $T=259120 349280 0 0 $X=258830 $Y=349045
X583 1 2 DCAP8BWP7T $T=263040 333600 1 0 $X=262750 $Y=329390
X584 1 2 DCAP8BWP7T $T=270880 302240 0 0 $X=270590 $Y=302005
X585 1 2 DCAP8BWP7T $T=273120 333600 1 0 $X=272830 $Y=329390
X586 1 2 DCAP8BWP7T $T=280960 357120 1 0 $X=280670 $Y=352910
X587 1 2 DCAP8BWP7T $T=287120 310080 1 0 $X=286830 $Y=305870
X588 1 2 DCAP8BWP7T $T=296640 341440 1 0 $X=296350 $Y=337230
X589 1 2 DCAP8BWP7T $T=300560 341440 0 0 $X=300270 $Y=341205
X590 1 2 DCAP8BWP7T $T=302240 333600 1 0 $X=301950 $Y=329390
X591 1 2 DCAP8BWP7T $T=307840 357120 1 0 $X=307550 $Y=352910
X592 1 2 DCAP8BWP7T $T=308960 317920 1 0 $X=308670 $Y=313710
X593 1 2 DCAP8BWP7T $T=310080 349280 1 0 $X=309790 $Y=345070
X594 1 2 DCAP8BWP7T $T=310640 325760 0 0 $X=310350 $Y=325525
X595 1 2 DCAP8BWP7T $T=320160 310080 1 0 $X=319870 $Y=305870
X596 1 2 DCAP8BWP7T $T=323520 302240 0 0 $X=323230 $Y=302005
X597 1 2 DCAP8BWP7T $T=323520 349280 0 0 $X=323230 $Y=349045
X598 1 2 DCAP8BWP7T $T=329120 341440 0 0 $X=328830 $Y=341205
X599 1 2 DCAP8BWP7T $T=342560 349280 0 0 $X=342270 $Y=349045
X600 1 2 DCAP8BWP7T $T=350960 325760 0 0 $X=350670 $Y=325525
X601 1 2 DCAP8BWP7T $T=364960 302240 1 0 $X=364670 $Y=298030
X602 1 2 DCAP8BWP7T $T=365520 325760 1 0 $X=365230 $Y=321550
X603 1 2 DCAP8BWP7T $T=365520 341440 1 0 $X=365230 $Y=337230
X604 1 2 DCAP8BWP7T $T=376160 310080 0 0 $X=375870 $Y=309845
X605 1 2 DCAP8BWP7T $T=389600 325760 1 0 $X=389310 $Y=321550
X606 1 2 DCAP8BWP7T $T=391840 325760 0 0 $X=391550 $Y=325525
X607 1 2 DCAP8BWP7T $T=395200 310080 1 0 $X=394910 $Y=305870
X608 1 2 DCAP8BWP7T $T=400800 325760 0 0 $X=400510 $Y=325525
X609 1 2 DCAP8BWP7T $T=404160 341440 1 0 $X=403870 $Y=337230
X610 1 2 DCAP8BWP7T $T=406960 310080 0 0 $X=406670 $Y=309845
X611 1 2 DCAP8BWP7T $T=422640 341440 0 0 $X=422350 $Y=341205
X612 1 2 DCAP8BWP7T $T=424320 333600 0 0 $X=424030 $Y=333365
X613 1 2 DCAP8BWP7T $T=433280 310080 0 0 $X=432990 $Y=309845
X614 1 2 DCAP8BWP7T $T=444480 341440 0 0 $X=444190 $Y=341205
X615 1 2 DCAP8BWP7T $T=446160 310080 0 0 $X=445870 $Y=309845
X616 1 2 DCAP8BWP7T $T=449520 357120 1 0 $X=449230 $Y=352910
X617 2 1 DCAPBWP7T $T=21120 333600 1 0 $X=20830 $Y=329390
X618 2 1 DCAPBWP7T $T=21120 349280 1 0 $X=20830 $Y=345070
X619 2 1 DCAPBWP7T $T=23360 341440 1 0 $X=23070 $Y=337230
X620 2 1 DCAPBWP7T $T=25040 294400 0 0 $X=24750 $Y=294165
X621 2 1 DCAPBWP7T $T=27280 333600 0 0 $X=26990 $Y=333365
X622 2 1 DCAPBWP7T $T=27840 349280 1 0 $X=27550 $Y=345070
X623 2 1 DCAPBWP7T $T=37360 333600 1 0 $X=37070 $Y=329390
X624 2 1 DCAPBWP7T $T=39600 294400 0 0 $X=39310 $Y=294165
X625 2 1 DCAPBWP7T $T=46320 302240 0 0 $X=46030 $Y=302005
X626 2 1 DCAPBWP7T $T=64240 349280 0 0 $X=63950 $Y=349045
X627 2 1 DCAPBWP7T $T=86640 310080 0 0 $X=86350 $Y=309845
X628 2 1 DCAPBWP7T $T=89440 333600 0 0 $X=89150 $Y=333365
X629 2 1 DCAPBWP7T $T=93920 341440 0 0 $X=93630 $Y=341205
X630 2 1 DCAPBWP7T $T=125840 349280 0 0 $X=125550 $Y=349045
X631 2 1 DCAPBWP7T $T=129760 349280 1 0 $X=129470 $Y=345070
X632 2 1 DCAPBWP7T $T=138160 302240 1 0 $X=137870 $Y=298030
X633 2 1 DCAPBWP7T $T=158320 310080 0 0 $X=158030 $Y=309845
X634 2 1 DCAPBWP7T $T=158320 317920 1 0 $X=158030 $Y=313710
X635 2 1 DCAPBWP7T $T=165600 325760 0 0 $X=165310 $Y=325525
X636 2 1 DCAPBWP7T $T=167840 349280 0 0 $X=167550 $Y=349045
X637 2 1 DCAPBWP7T $T=169520 310080 1 0 $X=169230 $Y=305870
X638 2 1 DCAPBWP7T $T=180160 302240 1 0 $X=179870 $Y=298030
X639 2 1 DCAPBWP7T $T=184080 310080 1 0 $X=183790 $Y=305870
X640 2 1 DCAPBWP7T $T=205360 302240 0 0 $X=205070 $Y=302005
X641 2 1 DCAPBWP7T $T=205360 310080 1 0 $X=205070 $Y=305870
X642 2 1 DCAPBWP7T $T=205360 349280 1 0 $X=205070 $Y=345070
X643 2 1 DCAPBWP7T $T=207600 317920 1 0 $X=207310 $Y=313710
X644 2 1 DCAPBWP7T $T=221040 349280 0 0 $X=220750 $Y=349045
X645 2 1 DCAPBWP7T $T=223840 302240 1 0 $X=223550 $Y=298030
X646 2 1 DCAPBWP7T $T=224400 302240 0 0 $X=224110 $Y=302005
X647 2 1 DCAPBWP7T $T=228320 333600 1 0 $X=228030 $Y=329390
X648 2 1 DCAPBWP7T $T=236720 341440 1 0 $X=236430 $Y=337230
X649 2 1 DCAPBWP7T $T=242320 325760 0 0 $X=242030 $Y=325525
X650 2 1 DCAPBWP7T $T=247360 302240 0 0 $X=247070 $Y=302005
X651 2 1 DCAPBWP7T $T=247360 325760 0 0 $X=247070 $Y=325525
X652 2 1 DCAPBWP7T $T=249600 341440 1 0 $X=249310 $Y=337230
X653 2 1 DCAPBWP7T $T=266960 349280 1 0 $X=266670 $Y=345070
X654 2 1 DCAPBWP7T $T=272000 302240 1 0 $X=271710 $Y=298030
X655 2 1 DCAPBWP7T $T=273680 349280 1 0 $X=273390 $Y=345070
X656 2 1 DCAPBWP7T $T=284320 317920 0 0 $X=284030 $Y=317685
X657 2 1 DCAPBWP7T $T=291600 325760 1 0 $X=291310 $Y=321550
X658 2 1 DCAPBWP7T $T=291600 333600 0 0 $X=291310 $Y=333365
X659 2 1 DCAPBWP7T $T=318480 294400 0 0 $X=318190 $Y=294165
X660 2 1 DCAPBWP7T $T=326320 325760 0 0 $X=326030 $Y=325525
X661 2 1 DCAPBWP7T $T=331360 349280 0 0 $X=331070 $Y=349045
X662 2 1 DCAPBWP7T $T=336960 325760 0 0 $X=336670 $Y=325525
X663 2 1 DCAPBWP7T $T=344800 349280 1 0 $X=344510 $Y=345070
X664 2 1 DCAPBWP7T $T=349280 341440 1 0 $X=348990 $Y=337230
X665 2 1 DCAPBWP7T $T=354320 317920 0 0 $X=354030 $Y=317685
X666 2 1 DCAPBWP7T $T=368320 294400 0 0 $X=368030 $Y=294165
X667 2 1 DCAPBWP7T $T=368320 325760 0 0 $X=368030 $Y=325525
X668 2 1 DCAPBWP7T $T=368320 333600 1 0 $X=368030 $Y=329390
X669 2 1 DCAPBWP7T $T=368320 349280 1 0 $X=368030 $Y=345070
X670 2 1 DCAPBWP7T $T=373360 294400 0 0 $X=373070 $Y=294165
X671 2 1 DCAPBWP7T $T=373360 341440 1 0 $X=373070 $Y=337230
X672 2 1 DCAPBWP7T $T=373360 349280 0 0 $X=373070 $Y=349045
X673 2 1 DCAPBWP7T $T=375600 349280 1 0 $X=375310 $Y=345070
X674 2 1 DCAPBWP7T $T=377840 310080 1 0 $X=377550 $Y=305870
X675 2 1 DCAPBWP7T $T=390720 294400 0 0 $X=390430 $Y=294165
X676 2 1 DCAPBWP7T $T=394640 310080 0 0 $X=394350 $Y=309845
X677 2 1 DCAPBWP7T $T=410320 325760 1 0 $X=410030 $Y=321550
X678 2 1 DCAPBWP7T $T=410320 349280 0 0 $X=410030 $Y=349045
X679 2 1 DCAPBWP7T $T=417600 302240 0 0 $X=417310 $Y=302005
X680 2 1 DCAPBWP7T $T=417600 349280 0 0 $X=417310 $Y=349045
X681 2 1 DCAPBWP7T $T=428800 302240 1 0 $X=428510 $Y=298030
X682 2 1 DCAPBWP7T $T=440560 341440 0 0 $X=440270 $Y=341205
X683 2 1 DCAPBWP7T $T=452320 302240 1 0 $X=452030 $Y=298030
X684 2 1 DCAPBWP7T $T=457360 357120 1 0 $X=457070 $Y=352910
X685 2 1 DCAPBWP7T $T=459600 310080 1 0 $X=459310 $Y=305870
X686 2 1 DCAPBWP7T $T=459600 317920 0 0 $X=459310 $Y=317685
X687 2 1 DCAPBWP7T $T=459600 341440 0 0 $X=459310 $Y=341205
X688 2 1 DCAPBWP7T $T=465200 333600 1 0 $X=464910 $Y=329390
X689 2 1 DCAPBWP7T $T=469120 317920 0 0 $X=468830 $Y=317685
X690 2 1 DCAPBWP7T $T=469120 349280 0 0 $X=468830 $Y=349045
X691 367 366 360 1175 1148 361 1 2 1171 AO222D0BWP7T $T=226640 317920 1 180 $X=220190 $Y=317685
X692 367 366 368 360 330 361 1 2 1161 AO222D0BWP7T $T=228320 325760 1 180 $X=221870 $Y=325525
X693 366 367 369 371 326 361 1 2 1177 AO222D0BWP7T $T=232240 302240 1 180 $X=225790 $Y=302005
X694 367 366 1175 365 325 361 1 2 1180 AO222D0BWP7T $T=226080 317920 1 0 $X=225790 $Y=313710
X695 366 367 373 374 375 361 1 2 1176 AO222D0BWP7T $T=228320 349280 1 0 $X=228030 $Y=345070
X696 366 367 374 364 376 361 1 2 1179 AO222D0BWP7T $T=236160 333600 0 180 $X=229710 $Y=329390
X697 366 367 383 373 384 361 1 2 388 AO222D0BWP7T $T=235040 357120 1 0 $X=234750 $Y=352910
X698 390 366 394 386 392 361 1 2 1183 AO222D0BWP7T $T=254080 333600 1 180 $X=247630 $Y=333365
X699 366 367 1192 1193 353 361 1 2 1189 AO222D0BWP7T $T=255200 341440 1 180 $X=248750 $Y=341205
X700 366 367 1195 387 396 361 1 2 1190 AO222D0BWP7T $T=256320 317920 0 180 $X=249870 $Y=313710
X701 366 367 401 1192 399 361 1 2 1191 AO222D0BWP7T $T=256880 325760 0 180 $X=250430 $Y=321550
X702 366 367 368 1205 402 361 1 2 1198 AO222D0BWP7T $T=259120 349280 1 180 $X=252670 $Y=349045
X703 366 367 409 1195 411 361 1 2 1211 AO222D0BWP7T $T=259680 317920 1 0 $X=259390 $Y=313710
X704 366 390 1193 386 412 361 1 2 1194 AO222D0BWP7T $T=259680 341440 0 0 $X=259390 $Y=341205
X705 539 367 1205 1294 546 361 1 2 1295 AO222D0BWP7T $T=353760 341440 0 0 $X=353470 $Y=341205
X706 539 367 1301 512 556 361 1 2 1306 AO222D0BWP7T $T=359920 349280 0 0 $X=359630 $Y=349045
X707 655 524 647 469 640 481 1 2 1349 AO222D0BWP7T $T=445040 310080 0 180 $X=438590 $Y=305870
X708 656 524 651 469 645 481 1 2 1351 AO222D0BWP7T $T=446160 310080 1 180 $X=439710 $Y=309845
X709 653 524 654 469 330 481 1 2 1327 AO222D0BWP7T $T=447280 302240 1 180 $X=440830 $Y=302005
X710 1354 524 660 469 1148 481 1 2 641 AO222D0BWP7T $T=447840 349280 0 180 $X=441390 $Y=345070
X711 662 524 659 469 652 481 1 2 644 AO222D0BWP7T $T=448400 341440 0 180 $X=441950 $Y=337230
X712 676 524 679 469 688 481 1 2 699 AO222D0BWP7T $T=462960 349280 0 0 $X=462670 $Y=349045
X713 665 1 384 1354 1358 2 1363 1364 OAI221D1BWP7T $T=460720 341440 1 0 $X=460430 $Y=337230
X714 1 2 ICV_4 $T=35120 341440 0 0 $X=34830 $Y=341205
X715 1 2 ICV_4 $T=54720 317920 1 0 $X=54430 $Y=313710
X716 1 2 ICV_4 $T=91680 333600 1 0 $X=91390 $Y=329390
X717 1 2 ICV_4 $T=102880 310080 0 0 $X=102590 $Y=309845
X718 1 2 ICV_4 $T=114080 349280 1 0 $X=113790 $Y=345070
X719 1 2 ICV_4 $T=209840 357120 1 0 $X=209550 $Y=352910
X720 1 2 ICV_4 $T=240080 310080 1 0 $X=239790 $Y=305870
X721 1 2 ICV_4 $T=240080 349280 1 0 $X=239790 $Y=345070
X722 1 2 ICV_4 $T=265840 341440 0 0 $X=265550 $Y=341205
X723 1 2 ICV_4 $T=282080 294400 0 0 $X=281790 $Y=294165
X724 1 2 ICV_4 $T=293280 294400 0 0 $X=292990 $Y=294165
X725 1 2 ICV_4 $T=300000 317920 1 0 $X=299710 $Y=313710
X726 1 2 ICV_4 $T=301680 325760 0 0 $X=301390 $Y=325525
X727 1 2 ICV_4 $T=324080 317920 0 0 $X=323790 $Y=317685
X728 1 2 ICV_4 $T=324080 333600 0 0 $X=323790 $Y=333365
X729 1 2 ICV_4 $T=343120 333600 1 0 $X=342830 $Y=329390
X730 1 2 ICV_4 $T=366080 349280 0 0 $X=365790 $Y=349045
X731 1 2 ICV_4 $T=408080 325760 0 0 $X=407790 $Y=325525
X732 1 2 ICV_4 $T=408080 349280 1 0 $X=407790 $Y=345070
X733 314 1132 303 2 1 298 DFCNQD1BWP7T $T=178480 341440 0 180 $X=165870 $Y=337230
X734 314 1133 303 2 1 1116 DFCNQD1BWP7T $T=178480 341440 1 180 $X=165870 $Y=341205
X735 314 1135 303 2 1 1119 DFCNQD1BWP7T $T=179600 325760 1 180 $X=166990 $Y=325525
X736 314 1137 303 2 1 1123 DFCNQD1BWP7T $T=181280 317920 0 180 $X=168670 $Y=313710
X737 314 1136 303 2 1 1124 DFCNQD1BWP7T $T=181280 333600 1 180 $X=168670 $Y=333365
X738 314 1144 303 2 1 1134 DFCNQD1BWP7T $T=188000 349280 1 180 $X=175390 $Y=349045
X739 314 1150 303 2 1 1141 DFCNQD1BWP7T $T=195280 341440 1 180 $X=182670 $Y=341205
X740 314 1152 303 2 1 1143 DFCNQD1BWP7T $T=196400 333600 1 180 $X=183790 $Y=333365
X741 314 1153 303 2 1 322 DFCNQD1BWP7T $T=196960 341440 0 180 $X=184350 $Y=337230
X742 314 1163 303 2 1 1145 DFCNQD1BWP7T $T=219360 302240 1 180 $X=206750 $Y=302005
X743 314 1165 303 2 1 1156 DFCNQD1BWP7T $T=221040 333600 1 180 $X=208430 $Y=333365
X744 314 1166 303 2 1 1149 DFCNQD1BWP7T $T=221040 341440 0 180 $X=208430 $Y=337230
X745 314 357 303 2 1 1157 DFCNQD1BWP7T $T=221040 349280 1 180 $X=208430 $Y=349045
X746 314 1167 303 2 1 1155 DFCNQD1BWP7T $T=221600 317920 0 180 $X=208990 $Y=313710
X747 314 1169 303 2 1 346 DFCNQD1BWP7T $T=223840 302240 0 180 $X=211230 $Y=298030
X748 314 1173 303 2 1 1151 DFCNQD1BWP7T $T=224400 310080 1 180 $X=211790 $Y=309845
X749 314 363 303 2 1 1147 DFCNQD1BWP7T $T=224960 341440 1 180 $X=212350 $Y=341205
X750 314 420 403 2 1 428 DFCNQD1BWP7T $T=266960 317920 1 0 $X=266670 $Y=313710
X751 530 526 523 2 1 508 DFCNQD1BWP7T $T=347040 302240 1 180 $X=334430 $Y=302005
X752 530 1327 523 2 1 1318 DFCNQD1BWP7T $T=404720 302240 1 180 $X=392110 $Y=302005
X753 530 1349 523 2 1 1350 DFCNQD1BWP7T $T=436080 325760 0 0 $X=435790 $Y=325525
X1066 1 2 ICV_8 $T=20000 333600 0 0 $X=19710 $Y=333365
X1067 1 2 ICV_8 $T=34000 349280 1 0 $X=33710 $Y=345070
X1068 1 2 ICV_8 $T=34000 357120 1 0 $X=33710 $Y=352910
X1069 1 2 ICV_8 $T=76000 333600 1 0 $X=75710 $Y=329390
X1070 1 2 ICV_8 $T=118000 333600 1 0 $X=117710 $Y=329390
X1071 1 2 ICV_8 $T=118000 341440 1 0 $X=117710 $Y=337230
X1072 1 2 ICV_8 $T=118000 349280 1 0 $X=117710 $Y=345070
X1073 1 2 ICV_8 $T=160000 302240 1 0 $X=159710 $Y=298030
X1074 1 2 ICV_8 $T=160000 302240 0 0 $X=159710 $Y=302005
X1075 1 2 ICV_8 $T=160000 310080 1 0 $X=159710 $Y=305870
X1076 1 2 ICV_8 $T=160000 310080 0 0 $X=159710 $Y=309845
X1077 1 2 ICV_8 $T=160000 317920 0 0 $X=159710 $Y=317685
X1078 1 2 ICV_8 $T=160000 325760 1 0 $X=159710 $Y=321550
X1079 1 2 ICV_8 $T=160000 333600 1 0 $X=159710 $Y=329390
X1080 1 2 ICV_8 $T=286000 317920 0 0 $X=285710 $Y=317685
X1081 1 2 ICV_8 $T=328000 317920 0 0 $X=327710 $Y=317685
X1082 1 2 ICV_8 $T=370000 310080 0 0 $X=369710 $Y=309845
X1083 1 2 ICV_8 $T=412000 317920 0 0 $X=411710 $Y=317685
X1084 1 2 ICV_8 $T=454000 333600 0 0 $X=453710 $Y=333365
X1085 1 2 ICV_8 $T=454000 341440 0 0 $X=453710 $Y=341205
X1086 1 2 ICV_9 $T=20000 325760 1 0 $X=19710 $Y=321550
X1087 1 2 ICV_9 $T=34000 294400 0 0 $X=33710 $Y=294165
X1088 1 2 ICV_9 $T=34000 310080 1 0 $X=33710 $Y=305870
X1089 1 2 ICV_9 $T=34000 310080 0 0 $X=33710 $Y=309845
X1090 1 2 ICV_9 $T=34000 317920 0 0 $X=33710 $Y=317685
X1091 1 2 ICV_9 $T=34000 325760 0 0 $X=33710 $Y=325525
X1092 1 2 ICV_9 $T=34000 333600 0 0 $X=33710 $Y=333365
X1093 1 2 ICV_9 $T=34000 349280 0 0 $X=33710 $Y=349045
X1094 1 2 ICV_9 $T=160000 317920 1 0 $X=159710 $Y=313710
X1095 1 2 ICV_9 $T=160000 325760 0 0 $X=159710 $Y=325525
X1096 1 2 ICV_9 $T=160000 333600 0 0 $X=159710 $Y=333365
X1097 1 2 ICV_9 $T=160000 341440 1 0 $X=159710 $Y=337230
X1098 1 2 ICV_9 $T=160000 341440 0 0 $X=159710 $Y=341205
X1099 1 2 ICV_9 $T=202000 294400 0 0 $X=201710 $Y=294165
X1100 1 2 ICV_9 $T=202000 302240 1 0 $X=201710 $Y=298030
X1101 1 2 ICV_9 $T=202000 317920 1 0 $X=201710 $Y=313710
X1102 1 2 ICV_9 $T=202000 333600 1 0 $X=201710 $Y=329390
X1103 1 2 ICV_9 $T=202000 333600 0 0 $X=201710 $Y=333365
X1104 1 2 ICV_9 $T=202000 349280 0 0 $X=201710 $Y=349045
X1105 1 2 ICV_9 $T=202000 357120 1 0 $X=201710 $Y=352910
X1106 1 2 ICV_9 $T=244000 310080 1 0 $X=243710 $Y=305870
X1107 1 2 ICV_9 $T=244000 310080 0 0 $X=243710 $Y=309845
X1108 1 2 ICV_9 $T=244000 317920 1 0 $X=243710 $Y=313710
X1109 1 2 ICV_9 $T=244000 325760 1 0 $X=243710 $Y=321550
X1110 1 2 ICV_9 $T=244000 341440 1 0 $X=243710 $Y=337230
X1111 1 2 ICV_9 $T=244000 349280 1 0 $X=243710 $Y=345070
X1112 1 2 ICV_9 $T=244000 349280 0 0 $X=243710 $Y=349045
X1113 1 2 ICV_9 $T=244000 357120 1 0 $X=243710 $Y=352910
X1114 1 2 ICV_9 $T=286000 325760 1 0 $X=285710 $Y=321550
X1115 1 2 ICV_9 $T=286000 333600 0 0 $X=285710 $Y=333365
X1116 1 2 ICV_9 $T=286000 341440 0 0 $X=285710 $Y=341205
X1117 1 2 ICV_9 $T=286000 349280 1 0 $X=285710 $Y=345070
X1118 1 2 ICV_9 $T=328000 302240 0 0 $X=327710 $Y=302005
X1119 1 2 ICV_9 $T=328000 310080 1 0 $X=327710 $Y=305870
X1120 1 2 ICV_9 $T=328000 317920 1 0 $X=327710 $Y=313710
X1121 1 2 ICV_9 $T=328000 325760 0 0 $X=327710 $Y=325525
X1122 1 2 ICV_9 $T=328000 333600 0 0 $X=327710 $Y=333365
X1123 1 2 ICV_9 $T=370000 317920 1 0 $X=369710 $Y=313710
X1124 1 2 ICV_9 $T=370000 325760 1 0 $X=369710 $Y=321550
X1125 1 2 ICV_9 $T=370000 333600 0 0 $X=369710 $Y=333365
X1126 1 2 ICV_9 $T=370000 349280 1 0 $X=369710 $Y=345070
X1127 1 2 ICV_9 $T=412000 294400 0 0 $X=411710 $Y=294165
X1128 1 2 ICV_9 $T=412000 302240 0 0 $X=411710 $Y=302005
X1129 1 2 ICV_9 $T=412000 325760 0 0 $X=411710 $Y=325525
X1130 1 2 ICV_9 $T=412000 341440 1 0 $X=411710 $Y=337230
X1131 1 2 ICV_9 $T=412000 349280 0 0 $X=411710 $Y=349045
X1132 1 2 ICV_9 $T=454000 302240 1 0 $X=453710 $Y=298030
X1133 1 2 ICV_9 $T=454000 302240 0 0 $X=453710 $Y=302005
X1134 1 2 ICV_9 $T=454000 310080 1 0 $X=453710 $Y=305870
X1135 1 2 ICV_9 $T=454000 310080 0 0 $X=453710 $Y=309845
X1136 1 2 ICV_9 $T=454000 317920 0 0 $X=453710 $Y=317685
X1137 1 2 ICV_9 $T=454000 325760 1 0 $X=453710 $Y=321550
X1138 1 2 ICV_9 $T=454000 325760 0 0 $X=453710 $Y=325525
X1139 1 2 ICV_9 $T=454000 333600 1 0 $X=453710 $Y=329390
X1140 1 2 ICV_9 $T=454000 341440 1 0 $X=453710 $Y=337230
X1141 1 2 ICV_10 $T=20000 294400 0 0 $X=19710 $Y=294165
X1142 1 2 ICV_10 $T=20000 317920 1 0 $X=19710 $Y=313710
X1143 1 2 ICV_10 $T=20000 341440 1 0 $X=19710 $Y=337230
X1144 1 2 ICV_10 $T=34000 333600 1 0 $X=33710 $Y=329390
X1145 1 2 ICV_10 $T=202000 302240 0 0 $X=201710 $Y=302005
X1146 1 2 ICV_10 $T=202000 310080 1 0 $X=201710 $Y=305870
X1147 1 2 ICV_10 $T=202000 349280 1 0 $X=201710 $Y=345070
X1148 1 2 ICV_10 $T=244000 302240 0 0 $X=243710 $Y=302005
X1149 1 2 ICV_10 $T=244000 325760 0 0 $X=243710 $Y=325525
X1150 1 2 ICV_10 $T=244000 341440 0 0 $X=243710 $Y=341205
X1151 1 2 ICV_10 $T=328000 349280 0 0 $X=327710 $Y=349045
X1152 1 2 ICV_10 $T=370000 294400 0 0 $X=369710 $Y=294165
X1153 1 2 ICV_10 $T=370000 325760 0 0 $X=369710 $Y=325525
X1154 1 2 ICV_10 $T=370000 341440 1 0 $X=369710 $Y=337230
X1155 1 2 ICV_10 $T=370000 349280 0 0 $X=369710 $Y=349045
X1156 1 2 ICV_10 $T=412000 333600 0 0 $X=411710 $Y=333365
X1157 1 2 ICV_10 $T=454000 357120 1 0 $X=453710 $Y=352910
X1189 1 2 ICV_13 $T=21120 310080 0 0 $X=20830 $Y=309845
X1190 1 2 ICV_13 $T=21120 317920 0 0 $X=20830 $Y=317685
X1191 1 2 ICV_13 $T=21120 325760 0 0 $X=20830 $Y=325525
X1192 1 2 ICV_13 $T=30640 310080 0 0 $X=30350 $Y=309845
X1193 1 2 ICV_13 $T=35120 302240 1 0 $X=34830 $Y=298030
X1194 1 2 ICV_13 $T=100640 294400 0 0 $X=100350 $Y=294165
X1195 1 2 ICV_13 $T=104560 325760 0 0 $X=104270 $Y=325525
X1196 1 2 ICV_13 $T=119120 310080 0 0 $X=118830 $Y=309845
X1197 1 2 ICV_13 $T=126960 302240 0 0 $X=126670 $Y=302005
X1198 1 2 ICV_13 $T=127520 333600 1 0 $X=127230 $Y=329390
X1199 1 2 ICV_13 $T=139280 317920 0 0 $X=138990 $Y=317685
X1200 1 2 ICV_13 $T=140400 325760 0 0 $X=140110 $Y=325525
X1201 1 2 ICV_13 $T=151040 325760 1 0 $X=150750 $Y=321550
X1202 1 2 ICV_13 $T=156640 310080 1 0 $X=156350 $Y=305870
X1203 1 2 ICV_13 $T=156640 317920 0 0 $X=156350 $Y=317685
X1204 1 2 ICV_13 $T=156640 341440 0 0 $X=156350 $Y=341205
X1205 1 2 ICV_13 $T=161120 349280 1 0 $X=160830 $Y=345070
X1206 1 2 ICV_13 $T=161120 357120 1 0 $X=160830 $Y=352910
X1207 1 2 ICV_13 $T=165600 317920 1 0 $X=165310 $Y=313710
X1208 1 2 ICV_13 $T=168960 349280 1 0 $X=168670 $Y=345070
X1209 1 2 ICV_13 $T=179600 333600 1 0 $X=179310 $Y=329390
X1210 1 2 ICV_13 $T=180720 357120 1 0 $X=180430 $Y=352910
X1211 1 2 ICV_13 $T=203120 310080 0 0 $X=202830 $Y=309845
X1212 1 2 ICV_13 $T=203120 317920 0 0 $X=202830 $Y=317685
X1213 1 2 ICV_13 $T=203120 325760 1 0 $X=202830 $Y=321550
X1214 1 2 ICV_13 $T=203120 325760 0 0 $X=202830 $Y=325525
X1215 1 2 ICV_13 $T=207600 333600 1 0 $X=207310 $Y=329390
X1216 1 2 ICV_13 $T=211520 325760 0 0 $X=211230 $Y=325525
X1217 1 2 ICV_13 $T=214320 310080 1 0 $X=214030 $Y=305870
X1218 1 2 ICV_13 $T=221040 357120 1 0 $X=220750 $Y=352910
X1219 1 2 ICV_13 $T=240640 302240 0 0 $X=240350 $Y=302005
X1220 1 2 ICV_13 $T=240640 325760 1 0 $X=240350 $Y=321550
X1221 1 2 ICV_13 $T=240640 341440 1 0 $X=240350 $Y=337230
X1222 1 2 ICV_13 $T=245120 317920 0 0 $X=244830 $Y=317685
X1223 1 2 ICV_13 $T=249600 349280 0 0 $X=249310 $Y=349045
X1224 1 2 ICV_13 $T=263600 349280 0 0 $X=263310 $Y=349045
X1225 1 2 ICV_13 $T=265840 317920 0 0 $X=265550 $Y=317685
X1226 1 2 ICV_13 $T=267520 333600 1 0 $X=267230 $Y=329390
X1227 1 2 ICV_13 $T=278160 302240 1 0 $X=277870 $Y=298030
X1228 1 2 ICV_13 $T=282640 310080 0 0 $X=282350 $Y=309845
X1229 1 2 ICV_13 $T=287120 294400 0 0 $X=286830 $Y=294165
X1230 1 2 ICV_13 $T=287120 325760 0 0 $X=286830 $Y=325525
X1231 1 2 ICV_13 $T=299440 325760 1 0 $X=299150 $Y=321550
X1232 1 2 ICV_13 $T=312320 357120 1 0 $X=312030 $Y=352910
X1233 1 2 ICV_13 $T=314560 349280 1 0 $X=314270 $Y=345070
X1234 1 2 ICV_13 $T=317360 317920 0 0 $X=317070 $Y=317685
X1235 1 2 ICV_13 $T=318480 357120 1 0 $X=318190 $Y=352910
X1236 1 2 ICV_13 $T=324640 310080 1 0 $X=324350 $Y=305870
X1237 1 2 ICV_13 $T=324640 357120 1 0 $X=324350 $Y=352910
X1238 1 2 ICV_13 $T=343120 325760 0 0 $X=342830 $Y=325525
X1239 1 2 ICV_13 $T=343680 341440 1 0 $X=343390 $Y=337230
X1240 1 2 ICV_13 $T=371120 317920 0 0 $X=370830 $Y=317685
X1241 1 2 ICV_13 $T=371120 333600 1 0 $X=370830 $Y=329390
X1242 1 2 ICV_13 $T=380080 357120 1 0 $X=379790 $Y=352910
X1243 1 2 ICV_13 $T=382320 302240 1 0 $X=382030 $Y=298030
X1244 1 2 ICV_13 $T=394080 325760 1 0 $X=393790 $Y=321550
X1245 1 2 ICV_13 $T=400800 349280 1 0 $X=400510 $Y=345070
X1246 1 2 ICV_13 $T=408640 341440 1 0 $X=408350 $Y=337230
X1247 1 2 ICV_13 $T=417600 294400 0 0 $X=417310 $Y=294165
X1248 1 2 ICV_13 $T=427120 341440 0 0 $X=426830 $Y=341205
X1249 1 2 ICV_13 $T=428800 333600 0 0 $X=428510 $Y=333365
X1250 1 2 ICV_13 $T=434400 349280 0 0 $X=434110 $Y=349045
X1251 1 2 ICV_13 $T=450640 310080 0 0 $X=450350 $Y=309845
X1252 1 2 ICV_13 $T=450640 333600 1 0 $X=450350 $Y=329390
X1253 1 2 ICV_13 $T=459600 333600 1 0 $X=459310 $Y=329390
X1254 1 2 ICV_13 $T=467440 325760 0 0 $X=467150 $Y=325525
X1255 305 301 2 301 1127 305 1 MAOI22D1BWP7T $T=177920 302240 0 180 $X=173150 $Y=298030
X1256 282 313 2 313 1138 282 1 MAOI22D1BWP7T $T=176240 317920 0 0 $X=175950 $Y=317685
X1257 277 321 2 321 1139 277 1 MAOI22D1BWP7T $T=193040 310080 1 180 $X=188270 $Y=309845
X1258 435 440 2 440 1223 435 1 MAOI22D1BWP7T $T=276480 357120 1 0 $X=276190 $Y=352910
X1259 410 1256 2 397 1263 499 1 MAOI22D1BWP7T $T=314560 341440 0 0 $X=314270 $Y=341205
X1260 497 500 2 500 1268 497 1 MAOI22D1BWP7T $T=324080 333600 1 180 $X=319310 $Y=333365
X1261 1275 520 2 520 1260 1275 1 MAOI22D1BWP7T $T=342560 349280 1 180 $X=337790 $Y=349045
X1262 1281 522 2 522 1266 1281 1 MAOI22D1BWP7T $T=343680 341440 0 180 $X=338910 $Y=337230
X1263 1314 566 2 566 572 1314 1 MAOI22D1BWP7T $T=377840 302240 1 0 $X=377550 $Y=298030
X1264 625 630 2 625 1289 630 1 MAOI22D1BWP7T $T=427680 317920 0 0 $X=427390 $Y=317685
X1265 1353 657 2 657 1345 1353 1 MAOI22D1BWP7T $T=448400 333600 1 180 $X=443630 $Y=333365
X1266 1357 666 2 664 1346 1357 1 MAOI22D1BWP7T $T=462400 333600 1 180 $X=457630 $Y=333365
X1267 8 1 2 13 INVD1BWP7T $T=23360 294400 0 0 $X=23070 $Y=294165
X1268 15 1 2 23 INVD1BWP7T $T=24480 310080 0 0 $X=24190 $Y=309845
X1269 31 1 2 24 INVD1BWP7T $T=28960 302240 1 180 $X=26990 $Y=302005
X1270 20 1 2 28 INVD1BWP7T $T=29520 333600 1 0 $X=29230 $Y=329390
X1271 38 1 2 870 INVD1BWP7T $T=31200 349280 0 180 $X=29230 $Y=345070
X1272 864 1 2 66 INVD1BWP7T $T=43520 317920 1 0 $X=43230 $Y=313710
X1273 77 1 2 876 INVD1BWP7T $T=49120 317920 0 180 $X=47150 $Y=313710
X1274 920 1 2 50 INVD1BWP7T $T=54160 341440 0 180 $X=52190 $Y=337230
X1275 934 1 2 169 INVD1BWP7T $T=86640 349280 1 0 $X=86350 $Y=345070
X1276 179 1 2 952 INVD1BWP7T $T=91120 294400 1 180 $X=89150 $Y=294165
X1277 172 1 2 967 INVD1BWP7T $T=92800 302240 1 0 $X=92510 $Y=298030
X1278 181 1 2 871 INVD1BWP7T $T=95040 349280 1 0 $X=94750 $Y=345070
X1279 226 1 2 885 INVD1BWP7T $T=114080 349280 0 180 $X=112110 $Y=345070
X1280 1065 1 2 212 INVD1BWP7T $T=129200 341440 0 180 $X=127230 $Y=337230
X1281 1037 1 2 240 INVD1BWP7T $T=140960 302240 0 0 $X=140670 $Y=302005
X1282 992 1 2 271 INVD1BWP7T $T=141520 294400 0 0 $X=141230 $Y=294165
X1283 257 1 2 274 INVD1BWP7T $T=153280 357120 0 180 $X=151310 $Y=352910
X1284 272 1 2 295 INVD1BWP7T $T=165600 325760 0 180 $X=163630 $Y=321550
X1285 1120 1 2 323 INVD1BWP7T $T=183520 294400 0 0 $X=183230 $Y=294165
X1286 576 1 2 1197 INVD1BWP7T $T=388480 310080 0 0 $X=388190 $Y=309845
X1287 1160 1 2 1321 INVD1BWP7T $T=395760 317920 1 0 $X=395470 $Y=313710
X1288 677 1 2 1314 INVD1BWP7T $T=464080 325760 0 180 $X=462110 $Y=321550
X1289 1 2 ICV_14 $T=42400 333600 1 0 $X=42110 $Y=329390
X1290 1 2 ICV_14 $T=154400 302240 1 0 $X=154110 $Y=298030
X1291 1 2 ICV_14 $T=196400 333600 1 0 $X=196110 $Y=329390
X1292 1 2 ICV_14 $T=196400 333600 0 0 $X=196110 $Y=333365
X1293 1 2 ICV_14 $T=196400 349280 1 0 $X=196110 $Y=345070
X1294 1 2 ICV_14 $T=196400 357120 1 0 $X=196110 $Y=352910
X1295 1 2 ICV_14 $T=203120 341440 1 0 $X=202830 $Y=337230
X1296 1 2 ICV_14 $T=221040 333600 0 0 $X=220750 $Y=333365
X1297 1 2 ICV_14 $T=221600 310080 1 0 $X=221310 $Y=305870
X1298 1 2 ICV_14 $T=238400 302240 1 0 $X=238110 $Y=298030
X1299 1 2 ICV_14 $T=280400 325760 0 0 $X=280110 $Y=325525
X1300 1 2 ICV_14 $T=280400 341440 1 0 $X=280110 $Y=337230
X1301 1 2 ICV_14 $T=280400 341440 0 0 $X=280110 $Y=341205
X1302 1 2 ICV_14 $T=280400 349280 1 0 $X=280110 $Y=345070
X1303 1 2 ICV_14 $T=315680 310080 0 0 $X=315390 $Y=309845
X1304 1 2 ICV_14 $T=339760 333600 0 0 $X=339470 $Y=333365
X1305 1 2 ICV_14 $T=345920 294400 0 0 $X=345630 $Y=294165
X1306 1 2 ICV_14 $T=349280 325760 1 0 $X=348990 $Y=321550
X1307 1 2 ICV_14 $T=378400 333600 0 0 $X=378110 $Y=333365
X1308 1 2 ICV_14 $T=386800 302240 0 0 $X=386510 $Y=302005
X1309 1 2 ICV_14 $T=389600 317920 0 0 $X=389310 $Y=317685
X1310 1 2 ICV_14 $T=390160 317920 1 0 $X=389870 $Y=313710
X1311 1 2 ICV_14 $T=406400 333600 0 0 $X=406110 $Y=333365
X1312 1 2 ICV_14 $T=422080 333600 1 0 $X=421790 $Y=329390
X1313 1 2 ICV_14 $T=448400 325760 0 0 $X=448110 $Y=325525
X1314 1 2 ICV_14 $T=448400 333600 0 0 $X=448110 $Y=333365
X1315 1 2 ICV_14 $T=455120 349280 0 0 $X=454830 $Y=349045
X1316 518 513 1 2 BUFFD2BWP7T $T=339760 317920 0 180 $X=336110 $Y=313710
X1317 675 667 1 2 BUFFD2BWP7T $T=463520 310080 1 180 $X=459870 $Y=309845
X1318 686 656 1 2 BUFFD2BWP7T $T=466320 310080 0 0 $X=466030 $Y=309845
X1319 705 695 1 2 BUFFD2BWP7T $T=470800 310080 0 180 $X=467150 $Y=305870
X1320 530 1351 523 633 1 2 DFCNQD2BWP7T $T=443360 302240 0 180 $X=430190 $Y=298030
X1321 1 2 DCAP16BWP7T $T=24480 341440 0 0 $X=24190 $Y=341205
X1322 1 2 DCAP16BWP7T $T=119120 294400 0 0 $X=118830 $Y=294165
X1323 1 2 DCAP16BWP7T $T=148240 325760 0 0 $X=147950 $Y=325525
X1324 1 2 DCAP16BWP7T $T=149360 317920 1 0 $X=149070 $Y=313710
X1325 1 2 DCAP16BWP7T $T=179600 349280 1 0 $X=179310 $Y=345070
X1326 1 2 DCAP16BWP7T $T=186880 302240 1 0 $X=186590 $Y=298030
X1327 1 2 DCAP16BWP7T $T=193040 310080 0 0 $X=192750 $Y=309845
X1328 1 2 DCAP16BWP7T $T=203120 341440 0 0 $X=202830 $Y=341205
X1329 1 2 DCAP16BWP7T $T=275920 325760 1 0 $X=275630 $Y=321550
X1330 1 2 DCAP16BWP7T $T=276480 310080 1 0 $X=276190 $Y=305870
X1331 1 2 DCAP16BWP7T $T=287120 349280 0 0 $X=286830 $Y=349045
X1332 1 2 DCAP16BWP7T $T=287120 357120 1 0 $X=286830 $Y=352910
X1333 1 2 DCAP16BWP7T $T=318480 302240 1 0 $X=318190 $Y=298030
X1334 1 2 DCAP16BWP7T $T=329120 294400 0 0 $X=328830 $Y=294165
X1335 1 2 DCAP16BWP7T $T=329120 302240 1 0 $X=328830 $Y=298030
X1336 1 2 DCAP16BWP7T $T=329120 341440 1 0 $X=328830 $Y=337230
X1337 1 2 DCAP16BWP7T $T=329120 349280 1 0 $X=328830 $Y=345070
X1338 1 2 DCAP16BWP7T $T=339760 310080 1 0 $X=339470 $Y=305870
X1339 1 2 DCAP16BWP7T $T=339760 317920 1 0 $X=339470 $Y=313710
X1340 1 2 DCAP16BWP7T $T=352640 333600 1 0 $X=352350 $Y=329390
X1341 1 2 DCAP16BWP7T $T=358240 357120 1 0 $X=357950 $Y=352910
X1342 1 2 DCAP16BWP7T $T=371120 341440 0 0 $X=370830 $Y=341205
X1343 1 2 DCAP16BWP7T $T=371120 357120 1 0 $X=370830 $Y=352910
X1344 1 2 DCAP16BWP7T $T=381200 317920 1 0 $X=380910 $Y=313710
X1345 1 2 DCAP16BWP7T $T=381760 294400 0 0 $X=381470 $Y=294165
X1346 1 2 DCAP16BWP7T $T=391840 349280 1 0 $X=391550 $Y=345070
X1347 1 2 DCAP16BWP7T $T=413120 349280 1 0 $X=412830 $Y=345070
X1348 1 2 DCAP16BWP7T $T=424320 310080 0 0 $X=424030 $Y=309845
X1349 1 2 DCAP16BWP7T $T=426000 357120 1 0 $X=425710 $Y=352910
X1350 1 2 DCAP16BWP7T $T=433840 294400 0 0 $X=433550 $Y=294165
X1351 1 2 DCAP16BWP7T $T=440000 317920 1 0 $X=439710 $Y=313710
X1352 1 2 DCAP16BWP7T $T=440560 357120 1 0 $X=440270 $Y=352910
X1353 1 2 DCAP16BWP7T $T=443360 302240 1 0 $X=443070 $Y=298030
X1354 1 2 DCAP16BWP7T $T=444480 349280 0 0 $X=444190 $Y=349045
X1355 863 1 2 5 CKND1BWP7T $T=21680 302240 0 0 $X=21390 $Y=302005
X1356 43 1 2 886 CKND1BWP7T $T=37920 349280 1 0 $X=37630 $Y=345070
X1357 58 1 2 51 CKND1BWP7T $T=43520 349280 0 180 $X=41550 $Y=345070
X1358 18 1 2 940 CKND1BWP7T $T=58640 325760 1 0 $X=58350 $Y=321550
X1359 173 1 2 27 CKND1BWP7T $T=87760 294400 0 0 $X=87470 $Y=294165
X1360 248 1 2 975 CKND1BWP7T $T=130320 310080 1 180 $X=128350 $Y=309845
X1361 284 1 2 1110 CKND1BWP7T $T=154400 302240 0 180 $X=152430 $Y=298030
X1362 265 1 2 290 CKND1BWP7T $T=156640 310080 0 180 $X=154670 $Y=305870
X1363 282 1 2 289 CKND1BWP7T $T=155520 294400 0 0 $X=155230 $Y=294165
X1364 370 366 1 2 INVD4BWP7T $T=228320 357120 0 180 $X=224110 $Y=352910
X1365 345 1 2 351 BUFFD3BWP7T $T=208720 294400 0 0 $X=208430 $Y=294165
X1366 356 1 2 1174 BUFFD3BWP7T $T=217680 310080 1 0 $X=217390 $Y=305870
X1367 516 1 2 524 BUFFD3BWP7T $T=338640 302240 1 0 $X=338350 $Y=298030
X1368 612 1 2 342 BUFFD3BWP7T $T=408080 349280 0 180 $X=403870 $Y=345070
X1369 707 1 2 689 BUFFD3BWP7T $T=470800 325760 0 180 $X=466590 $Y=321550
X1370 690 1 2 696 BUFFD3BWP7T $T=466880 333600 1 0 $X=466590 $Y=329390
X1371 1154 328 320 1 2 CKXOR2D4BWP7T $T=196400 357120 0 180 $X=183790 $Y=352910
X1372 1265 484 472 1 2 CKXOR2D4BWP7T $T=317360 317920 1 180 $X=304750 $Y=317685
X1373 212 1033 2 973 1 198 1034 AOI22D1BWP7T $T=106240 325760 0 180 $X=102030 $Y=321550
X1374 282 1110 2 289 1 284 287 AOI22D1BWP7T $T=155520 294400 1 180 $X=151310 $Y=294165
X1375 277 1114 2 297 1 1112 1121 AOI22D1BWP7T $T=167840 310080 1 180 $X=163630 $Y=309845
X1376 1114 295 2 1112 1 272 1118 AOI22D1BWP7T $T=163920 317920 0 0 $X=163630 $Y=317685
X1377 400 391 2 1199 1 397 406 AOI22D1BWP7T $T=254080 302240 0 0 $X=253790 $Y=302005
X1378 398 1207 2 395 1 1185 1210 AOI22D1BWP7T $T=259120 302240 0 0 $X=258830 $Y=302005
X1379 481 479 2 469 1 476 1225 AOI22D1BWP7T $T=310080 349280 0 180 $X=305870 $Y=345070
X1380 398 1259 2 395 1 1255 1261 AOI22D1BWP7T $T=308400 333600 1 0 $X=308110 $Y=329390
X1381 481 494 2 469 1 486 1262 AOI22D1BWP7T $T=319040 325760 1 180 $X=314830 $Y=325525
X1382 481 342 2 469 1 1216 496 AOI22D1BWP7T $T=321840 349280 0 180 $X=317630 $Y=345070
X1383 481 502 2 469 1 491 1269 AOI22D1BWP7T $T=325200 341440 1 180 $X=320990 $Y=341205
X1384 1303 547 2 1299 1 552 1309 AOI22D1BWP7T $T=373920 302240 0 0 $X=373630 $Y=302005
X1385 481 578 2 469 1 575 1316 AOI22D1BWP7T $T=386800 325760 1 180 $X=382590 $Y=325525
X1386 1324 1160 2 1294 1 1321 596 AOI22D1BWP7T $T=396320 333600 0 0 $X=396030 $Y=333365
X1387 1338 1174 2 1339 1 1321 1331 AOI22D1BWP7T $T=420400 310080 0 0 $X=420110 $Y=309845
X1388 439 1224 2 446 1152 1 OAI21D1BWP7T $T=277040 341440 1 0 $X=276750 $Y=337230
X1389 452 448 2 1231 1226 1 OAI21D1BWP7T $T=293280 333600 0 180 $X=289630 $Y=329390
X1390 408 1270 2 1252 1271 1 OAI21D1BWP7T $T=324080 317920 1 180 $X=320430 $Y=317685
X1391 408 1272 2 1273 1265 1 OAI21D1BWP7T $T=320720 325760 0 0 $X=320430 $Y=325525
X1392 551 1345 2 636 1307 1 OAI21D1BWP7T $T=423760 310080 1 0 $X=423470 $Y=305870
X1393 551 1346 2 631 1283 1 OAI21D1BWP7T $T=427680 333600 1 0 $X=427390 $Y=329390
X1394 635 1332 2 1348 1330 1 OAI21D1BWP7T $T=433840 341440 1 180 $X=430190 $Y=341205
X1395 408 1352 2 1343 639 1 OAI21D1BWP7T $T=440000 325760 1 0 $X=439710 $Y=321550
X1396 339 2 314 1 CKND12BWP7T $T=206480 317920 0 0 $X=206190 $Y=317685
X1397 336 303 1 2 BUFFD6BWP7T $T=196400 349280 0 180 $X=189390 $Y=345070
X1398 865 4 2 1 INVD2BWP7T $T=23360 349280 1 180 $X=20830 $Y=349045
X1399 10 6 2 1 INVD2BWP7T $T=24480 341440 1 180 $X=21950 $Y=341205
X1400 877 35 2 1 INVD2BWP7T $T=31200 333600 1 180 $X=28670 $Y=333365
X1401 84 93 2 1 INVD2BWP7T $T=54160 357120 0 180 $X=51630 $Y=352910
X1402 268 267 2 1 INVD2BWP7T $T=153280 349280 0 180 $X=150750 $Y=345070
X1403 1131 352 2 1 INVD2BWP7T $T=212080 310080 1 0 $X=211790 $Y=305870
X1404 445 423 2 1 INVD2BWP7T $T=279840 294400 0 0 $X=279550 $Y=294165
X1405 550 557 2 1 INVD2BWP7T $T=363280 325760 1 0 $X=362990 $Y=321550
X1406 484 559 2 1 INVD2BWP7T $T=376160 310080 1 180 $X=373630 $Y=309845
X1407 578 553 2 1 INVD2BWP7T $T=385120 317920 0 0 $X=384830 $Y=317685
X1408 593 595 2 1 INVD2BWP7T $T=396320 310080 0 0 $X=396030 $Y=309845
X1409 597 610 2 1 INVD2BWP7T $T=432160 333600 0 0 $X=431870 $Y=333365
X1410 646 634 2 1 INVD2BWP7T $T=442240 341440 0 0 $X=441950 $Y=341205
X1411 293 301 1 2 1126 CKXOR2D1BWP7T $T=166160 302240 1 0 $X=165870 $Y=298030
X1412 318 317 1 2 1142 CKXOR2D1BWP7T $T=181840 302240 1 0 $X=181550 $Y=298030
X1413 1159 342 1 2 1098 CKXOR2D1BWP7T $T=211520 325760 1 180 $X=206190 $Y=325525
X1414 1175 377 1 2 1181 CKXOR2D1BWP7T $T=229440 317920 0 0 $X=229150 $Y=317685
X1415 377 383 1 2 1188 CKXOR2D1BWP7T $T=235040 325760 0 0 $X=234750 $Y=325525
X1416 1184 382 1 2 1109 CKXOR2D1BWP7T $T=240080 349280 0 180 $X=234750 $Y=345070
X1417 389 393 1 2 1196 CKXOR2D1BWP7T $T=247920 294400 0 0 $X=247630 $Y=294165
X1418 391 1195 1 2 1199 CKXOR2D1BWP7T $T=249040 302240 0 0 $X=248750 $Y=302005
X1419 422 424 1 2 1221 CKXOR2D1BWP7T $T=269760 341440 0 0 $X=269470 $Y=341205
X1420 478 486 1 2 1254 CKXOR2D1BWP7T $T=308960 294400 0 0 $X=308670 $Y=294165
X1421 1187 487 1 2 1257 CKXOR2D1BWP7T $T=310640 310080 0 0 $X=310350 $Y=309845
X1422 1267 491 1 2 1264 CKXOR2D1BWP7T $T=320160 310080 0 180 $X=314830 $Y=305870
X1423 1304 554 1 2 1300 CKXOR2D1BWP7T $T=365520 341440 0 180 $X=360190 $Y=337230
X1424 1322 602 1 2 1329 CKXOR2D1BWP7T $T=398560 349280 0 0 $X=398270 $Y=349045
X1425 622 1321 1 2 1344 CKXOR2D1BWP7T $T=422080 317920 1 0 $X=421790 $Y=313710
X1426 1164 353 350 1 2 CKXOR2D2BWP7T $T=218800 325760 0 180 $X=212350 $Y=321550
X1427 441 428 279 1 2 CKXOR2D2BWP7T $T=279280 310080 1 180 $X=272830 $Y=309845
X1428 1237 459 1102 1 2 CKXOR2D2BWP7T $T=300560 341440 1 180 $X=294110 $Y=341205
X1429 1271 495 489 1 2 CKXOR2D2BWP7T $T=323520 302240 1 180 $X=317070 $Y=302005
X1430 517 509 296 1 2 CKXOR2D2BWP7T $T=339760 310080 0 180 $X=333310 $Y=305870
X1431 1285 528 1108 1 2 CKXOR2D2BWP7T $T=349280 325760 0 180 $X=342830 $Y=321550
X1432 603 597 269 1 2 CKXOR2D2BWP7T $T=403600 325760 0 180 $X=397150 $Y=321550
X1433 2 1 DCAP32BWP7T $T=224960 341440 0 0 $X=224670 $Y=341205
X1434 2 1 DCAP32BWP7T $T=305600 349280 0 0 $X=305310 $Y=349045
X1435 2 1 DCAP32BWP7T $T=310080 325760 1 0 $X=309790 $Y=321550
X1436 1139 1134 1131 1127 290 1 2 XNR4D1BWP7T $T=184080 310080 0 180 $X=170910 $Y=305870
X1437 362 1 2 353 BUFFD5BWP7T $T=222160 349280 0 180 $X=215710 $Y=345070
X1438 1232 1233 454 398 1 2 OAI21D0BWP7T $T=290480 294400 0 0 $X=290190 $Y=294165
X1439 455 1242 457 426 1 2 OAI21D0BWP7T $T=297200 310080 1 0 $X=296910 $Y=305870
X1440 1241 1246 462 426 1 2 OAI21D0BWP7T $T=298880 325760 0 0 $X=298590 $Y=325525
X1441 464 1250 470 398 1 2 OAI21D0BWP7T $T=302800 310080 1 0 $X=302510 $Y=305870
X1442 507 1276 515 1280 1 2 OAI21D0BWP7T $T=336960 341440 0 0 $X=336670 $Y=341205
X1443 1286 1290 535 398 1 2 OAI21D0BWP7T $T=350960 341440 1 0 $X=350670 $Y=337230
X1444 1305 1317 563 426 1 2 OAI21D0BWP7T $T=375040 341440 1 0 $X=374750 $Y=337230
X1445 1309 1319 573 398 1 2 OAI21D0BWP7T $T=381760 341440 1 0 $X=381470 $Y=337230
X1446 614 1340 617 1347 1 2 OAI21D0BWP7T $T=417600 325760 0 0 $X=417310 $Y=325525
X1447 1333 1341 623 398 1 2 OAI21D0BWP7T $T=421520 333600 0 0 $X=421230 $Y=333365
X1448 1121 1123 310 311 317 1 2 XNR4D0BWP7T $T=168400 294400 0 0 $X=168110 $Y=294165
X1449 1116 1118 312 315 294 1 2 XNR4D0BWP7T $T=168960 310080 0 0 $X=168670 $Y=309845
X1450 1141 1138 1128 1127 272 1 2 XNR4D0BWP7T $T=182960 325760 0 180 $X=169790 $Y=321550
X1451 1125 1145 1140 1139 316 1 2 XNR4D0BWP7T $T=190240 302240 1 180 $X=177070 $Y=302005
X1452 1125 1143 325 1138 319 1 2 XNR4D2BWP7T $T=195280 317920 1 180 $X=181550 $Y=317685
X1453 329 1149 326 282 1142 1 2 XNR4D2BWP7T $T=196400 333600 0 180 $X=182670 $Y=329390
X1454 1130 1151 327 1146 321 1 2 XNR4D2BWP7T $T=197520 317920 0 180 $X=183790 $Y=313710
X1455 1126 1147 334 286 337 1 2 XNR4D2BWP7T $T=185760 294400 0 0 $X=185470 $Y=294165
X1456 338 1155 330 1126 324 1 2 XNR4D2BWP7T $T=199200 310080 0 180 $X=185470 $Y=305870
X1457 277 1156 1148 1146 1142 1 2 XNR4D2BWP7T $T=199200 325760 0 180 $X=185470 $Y=321550
X1458 1130 1157 331 329 313 1 2 XNR4D2BWP7T $T=199200 325760 1 180 $X=185470 $Y=325525
X1459 1114 1119 1112 1 2 307 MUX2ND1BWP7T $T=169520 317920 0 0 $X=169230 $Y=317685
X1460 1118 292 1 2 1130 XNR2D1BWP7T $T=170640 302240 0 0 $X=170350 $Y=302005
X1461 371 385 1 2 1185 XNR2D1BWP7T $T=235600 302240 0 0 $X=235310 $Y=302005
X1462 369 344 1 2 1187 XNR2D1BWP7T $T=235600 317920 1 0 $X=235310 $Y=313710
X1463 1181 1197 1 2 1201 XNR2D1BWP7T $T=249600 310080 0 0 $X=249310 $Y=309845
X1464 1202 1192 1 2 1206 XNR2D1BWP7T $T=254640 333600 0 0 $X=254350 $Y=333365
X1465 1185 419 1 2 1207 XNR2D1BWP7T $T=265840 302240 0 0 $X=265550 $Y=302005
X1466 1193 347 1 2 1220 XNR2D1BWP7T $T=268640 349280 1 0 $X=268350 $Y=345070
X1467 463 467 1 2 1249 XNR2D1BWP7T $T=297200 294400 0 0 $X=296910 $Y=294165
X1468 1205 473 1 2 1255 XNR2D1BWP7T $T=304480 341440 1 0 $X=304190 $Y=337230
X1469 1255 480 1 2 1259 XNR2D1BWP7T $T=305600 325760 0 0 $X=305310 $Y=325525
X1470 504 445 1 2 1267 XNR2D1BWP7T $T=325200 294400 1 180 $X=319870 $Y=294165
X1471 1256 512 1 2 499 XNR2D1BWP7T $T=333040 349280 0 0 $X=332750 $Y=349045
X1472 545 550 1 2 1304 XNR2D1BWP7T $T=356560 333600 0 0 $X=356270 $Y=333365
X1473 582 586 1 2 1322 XNR2D1BWP7T $T=386240 349280 0 0 $X=385950 $Y=349045
X1474 502 587 2 1 CKND2BWP7T $T=389600 325760 0 0 $X=389310 $Y=325525
X1475 494 607 2 1 CKND2BWP7T $T=403040 317920 0 0 $X=402750 $Y=317685
X1476 7 1 2 3 CKND0BWP7T $T=23360 357120 0 180 $X=21390 $Y=352910
X1477 64 1 2 1027 CKND0BWP7T $T=101200 341440 1 0 $X=100910 $Y=337230
X1478 917 1 2 198 CKND0BWP7T $T=104560 325760 1 180 $X=102590 $Y=325525
X1479 1108 1 2 1099 CKND0BWP7T $T=151040 310080 1 180 $X=149070 $Y=309845
X1480 265 2 1110 292 284 290 1 AOI22D2BWP7T $T=150480 302240 0 0 $X=150190 $Y=302005
X1481 293 2 1113 1125 294 1117 1 AOI22D2BWP7T $T=163920 302240 0 0 $X=163630 $Y=302005
X1482 381 2 378 1186 380 387 1 AOI22D2BWP7T $T=234480 317920 0 0 $X=234190 $Y=317685
X1483 521 2 445 1278 423 525 1 AOI22D2BWP7T $T=339200 294400 0 0 $X=338910 $Y=294165
X1484 481 2 484 540 1282 469 1 AOI22D2BWP7T $T=347040 349280 0 0 $X=346750 $Y=349045
X1485 1292 2 547 1298 552 1297 1 AOI22D2BWP7T $T=356000 317920 0 0 $X=355710 $Y=317685
X1486 568 2 547 1293 552 561 1 AOI22D2BWP7T $T=381760 294400 1 180 $X=374750 $Y=294165
X1487 481 2 546 571 574 469 1 AOI22D2BWP7T $T=387360 310080 1 180 $X=380350 $Y=309845
X1488 481 2 588 1248 576 469 1 AOI22D2BWP7T $T=389600 325760 0 180 $X=382590 $Y=321550
X1489 1301 2 1160 589 1321 584 1 AOI22D2BWP7T $T=384000 333600 0 0 $X=383710 $Y=333365
X1490 481 2 569 579 581 469 1 AOI22D2BWP7T $T=392400 302240 0 180 $X=385390 $Y=298030
X1491 1328 2 1174 1332 1321 604 1 AOI22D2BWP7T $T=401360 310080 1 0 $X=401070 $Y=305870
X1492 481 2 638 650 649 469 1 AOI22D2BWP7T $T=437760 349280 0 0 $X=437470 $Y=349045
X1493 1124 1129 1115 308 1 2 MUX2ND0BWP7T $T=179600 333600 0 180 $X=174830 $Y=329390
X1494 1188 1216 1218 1219 1 2 MUX2ND0BWP7T $T=269200 317920 0 0 $X=268910 $Y=317685
X1495 1199 425 431 427 1 2 MUX2ND0BWP7T $T=272000 310080 1 0 $X=271710 $Y=305870
X1496 1196 430 436 1209 1 2 MUX2ND0BWP7T $T=273680 302240 1 0 $X=273390 $Y=298030
X1497 1206 432 438 1213 1 2 MUX2ND0BWP7T $T=274240 333600 0 0 $X=273950 $Y=333365
X1498 1221 443 435 1215 1 2 MUX2ND0BWP7T $T=280400 341440 1 180 $X=275630 $Y=341205
X1499 1220 468 466 1247 1 2 MUX2ND0BWP7T $T=302800 357120 0 180 $X=298030 $Y=352910
X1500 1249 505 1275 1270 1 2 MUX2ND0BWP7T $T=336400 317920 1 180 $X=331630 $Y=317685
X1501 510 1282 1281 1272 1 2 MUX2ND0BWP7T $T=343120 325760 1 180 $X=338350 $Y=325525
X1502 1293 562 1313 1311 1 2 MUX2ND0BWP7T $T=374480 317920 0 0 $X=374190 $Y=317685
X1503 1344 649 1353 1352 1 2 MUX2ND0BWP7T $T=442800 317920 0 0 $X=442510 $Y=317685
X1504 1038 1044 1045 212 1028 2 1 AOI22D0BWP7T $T=112400 325760 0 180 $X=108750 $Y=321550
X1505 1201 1200 1181 398 395 2 1 AOI22D0BWP7T $T=255760 310080 0 180 $X=252110 $Y=305870
X1506 400 1203 1196 393 397 2 1 AOI22D0BWP7T $T=256320 294400 1 180 $X=252670 $Y=294165
X1507 377 1204 397 400 1188 2 1 AOI22D0BWP7T $T=255760 310080 0 0 $X=255470 $Y=309845
X1508 210 1 2 1059 CKBD0BWP7T $T=121920 333600 1 0 $X=121630 $Y=329390
X1509 348 1 2 1154 CKBD0BWP7T $T=209840 357120 0 180 $X=207310 $Y=352910
X1510 385 1 2 1202 CKBD0BWP7T $T=238960 333600 1 0 $X=238670 $Y=329390
X1511 429 1 2 1222 CKBD0BWP7T $T=274240 294400 0 0 $X=273950 $Y=294165
X1512 473 1 2 1256 CKBD0BWP7T $T=305040 341440 0 0 $X=304750 $Y=341205
X1513 669 1 2 666 CKBD0BWP7T $T=462400 325760 0 180 $X=459870 $Y=321550
X1514 41 2 889 890 1 NR2D1BWP7T $T=39600 310080 0 0 $X=39310 $Y=309845
X1515 65 2 893 887 1 NR2D1BWP7T $T=45760 349280 0 180 $X=43230 $Y=345070
X1516 58 2 899 887 1 NR2D1BWP7T $T=46320 341440 1 180 $X=43790 $Y=341205
X1517 78 2 898 890 1 NR2D1BWP7T $T=50240 302240 1 180 $X=47710 $Y=302005
X1518 966 2 972 977 1 NR2D1BWP7T $T=70960 325760 0 0 $X=70670 $Y=325525
X1519 967 2 990 176 1 NR2D1BWP7T $T=91680 310080 0 180 $X=89150 $Y=305870
X1520 186 2 174 950 1 NR2D1BWP7T $T=93360 333600 1 180 $X=90830 $Y=333365
X1521 921 2 1049 215 1 NR2D1BWP7T $T=112400 341440 0 0 $X=112110 $Y=341205
X1522 264 2 283 285 1 NR2D1BWP7T $T=148240 357120 1 0 $X=147950 $Y=352910
X1523 467 2 1234 421 1 NR2D1BWP7T $T=302800 302240 0 180 $X=300270 $Y=298030
X1524 1000 1048 212 1063 1 2 AOI21D0BWP7T $T=123040 325760 1 0 $X=122750 $Y=321550
X1525 1029 1062 240 1050 1 2 AOI21D0BWP7T $T=124160 302240 0 0 $X=123870 $Y=302005
X1526 448 1231 452 408 1 2 AOI21D0BWP7T $T=290480 325760 0 0 $X=290190 $Y=325525
X1527 1232 1230 454 1233 1 2 AOI21D0BWP7T $T=292720 302240 1 0 $X=292430 $Y=298030
X1528 455 1236 457 1242 1 2 AOI21D0BWP7T $T=293280 310080 1 0 $X=292990 $Y=305870
X1529 1241 1244 462 1246 1 2 AOI21D0BWP7T $T=296080 325760 0 0 $X=295790 $Y=325525
X1530 1247 1235 426 1251 1 2 AOI21D0BWP7T $T=300000 349280 1 0 $X=299710 $Y=345070
X1531 464 1245 470 1250 1 2 AOI21D0BWP7T $T=301120 310080 0 0 $X=300830 $Y=309845
X1532 507 1280 515 408 1 2 AOI21D0BWP7T $T=336960 333600 0 0 $X=336670 $Y=333365
X1533 1311 1296 426 560 1 2 AOI21D0BWP7T $T=377840 325760 1 180 $X=374750 $Y=325525
X1534 1305 1310 563 1317 1 2 AOI21D0BWP7T $T=375600 333600 0 0 $X=375310 $Y=333365
X1535 1309 1312 573 1319 1 2 AOI21D0BWP7T $T=380080 333600 1 0 $X=379790 $Y=329390
X1536 1333 1342 623 1341 1 2 AOI21D0BWP7T $T=422080 341440 1 0 $X=421790 $Y=337230
X1537 614 1347 617 408 1 2 AOI21D0BWP7T $T=429920 325760 1 0 $X=429630 $Y=321550
X1538 1332 1348 635 408 1 2 AOI21D0BWP7T $T=432160 341440 1 0 $X=431870 $Y=337230
X1539 878 875 23 24 2 1 18 NR4D1BWP7T $T=30640 310080 0 180 $X=24750 $Y=305870
X1540 880 34 28 870 2 1 21 NR4D1BWP7T $T=30640 341440 0 180 $X=24750 $Y=337230
X1541 881 32 863 25 2 1 867 NR4D1BWP7T $T=31200 317920 0 180 $X=25310 $Y=313710
X1542 897 864 24 884 2 1 41 NR4D1BWP7T $T=44080 302240 0 180 $X=38190 $Y=298030
X1543 895 906 87 74 2 1 883 NR4D1BWP7T $T=52480 349280 0 180 $X=46590 $Y=345070
X1544 918 89 35 910 2 1 76 NR4D1BWP7T $T=53600 333600 0 180 $X=47710 $Y=329390
X1545 922 876 94 82 2 1 868 NR4D1BWP7T $T=54720 317920 0 180 $X=48830 $Y=313710
X1546 912 89 931 937 2 1 942 NR4D1BWP7T $T=55280 333600 1 0 $X=54990 $Y=329390
X1547 955 126 870 118 2 1 58 NR4D1BWP7T $T=65920 349280 0 180 $X=60030 $Y=345070
X1548 978 144 135 904 2 1 116 NR4D1BWP7T $T=73200 302240 0 180 $X=67310 $Y=298030
X1549 147 141 93 921 2 1 65 NR4D1BWP7T $T=73200 357120 0 180 $X=67310 $Y=352910
X1550 970 159 158 979 2 1 130 NR4D1BWP7T $T=85520 294400 1 180 $X=79630 $Y=294165
X1551 993 874 160 148 2 1 949 NR4D1BWP7T $T=86640 325760 1 180 $X=80750 $Y=325525
X1552 924 138 982 154 2 1 152 NR4D1BWP7T $T=87200 310080 0 180 $X=81310 $Y=305870
X1553 178 100 195 200 2 1 936 NR4D1BWP7T $T=93920 317920 0 0 $X=93630 $Y=317685
X1554 1024 971 1007 1011 2 1 186 NR4D1BWP7T $T=101200 333600 0 180 $X=95310 $Y=329390
X1555 1039 216 214 939 2 1 211 NR4D1BWP7T $T=109600 294400 1 180 $X=103710 $Y=294165
X1556 1047 214 218 213 2 1 144 NR4D1BWP7T $T=111280 302240 1 180 $X=105390 $Y=302005
X1557 1055 949 215 222 2 1 227 NR4D1BWP7T $T=114080 357120 0 180 $X=108190 $Y=352910
X1558 1061 89 219 994 2 1 1066 NR4D1BWP7T $T=121920 341440 1 0 $X=121630 $Y=337230
X1559 917 2 933 97 912 96 1 AOI31D2BWP7T $T=51920 325760 0 0 $X=51630 $Y=325525
X1560 170 2 947 269 79 267 1 AOI31D2BWP7T $T=139280 341440 0 0 $X=138990 $Y=341205
X1561 21 906 907 911 1 2 914 OA31D0BWP7T $T=45760 333600 0 0 $X=45470 $Y=333365
X1562 930 114 941 911 1 2 945 OA31D0BWP7T $T=58640 325760 0 0 $X=58350 $Y=325525
X1563 249 959 1071 1045 1 2 1083 OA31D0BWP7T $T=130880 333600 1 0 $X=130590 $Y=329390
X1564 268 269 273 226 1 2 1111 OA31D0BWP7T $T=156640 341440 1 180 $X=151870 $Y=341205
X1565 9 1 868 17 2 ND2D1BWP7T $T=23360 317920 1 0 $X=23070 $Y=313710
X1566 6 1 12 7 2 ND2D1BWP7T $T=25600 357120 0 180 $X=23070 $Y=352910
X1567 4 1 30 26 2 ND2D1BWP7T $T=27280 357120 1 0 $X=26990 $Y=352910
X1568 31 1 37 29 2 ND2D1BWP7T $T=28960 302240 0 0 $X=28670 $Y=302005
X1569 6 1 877 39 2 ND2D1BWP7T $T=28960 349280 0 0 $X=28670 $Y=349045
X1570 44 1 883 30 2 ND2D1BWP7T $T=40160 357120 0 180 $X=37630 $Y=352910
X1571 56 1 884 45 2 ND2D1BWP7T $T=43520 294400 1 180 $X=40990 $Y=294165
X1572 67 1 63 54 2 ND2D1BWP7T $T=46320 302240 0 180 $X=43790 $Y=298030
X1573 79 1 84 39 2 ND2D1BWP7T $T=49120 357120 1 0 $X=48830 $Y=352910
X1574 51 1 910 103 2 ND2D1BWP7T $T=53600 349280 1 0 $X=53310 $Y=345070
X1575 110 1 101 26 2 ND2D1BWP7T $T=58080 357120 0 180 $X=55550 $Y=352910
X1576 40 1 932 113 2 ND2D1BWP7T $T=56960 302240 0 0 $X=56670 $Y=302005
X1577 109 1 118 873 2 ND2D1BWP7T $T=57520 341440 0 0 $X=57230 $Y=341205
X1578 110 1 934 69 2 ND2D1BWP7T $T=60320 357120 0 180 $X=57790 $Y=352910
X1579 932 1 936 940 2 ND2D1BWP7T $T=58640 317920 1 0 $X=58350 $Y=313710
X1580 871 1 958 101 2 ND2D1BWP7T $T=70400 349280 0 180 $X=67870 $Y=345070
X1581 129 1 971 964 2 ND2D1BWP7T $T=73200 333600 0 180 $X=70670 $Y=329390
X1582 150 1 981 934 2 ND2D1BWP7T $T=82160 349280 0 180 $X=79630 $Y=345070
X1583 940 1 167 986 2 ND2D1BWP7T $T=85520 294400 0 0 $X=85230 $Y=294165
X1584 197 1 1007 1018 2 ND2D1BWP7T $T=96720 349280 0 0 $X=96430 $Y=349045
X1585 6 1 120 201 2 ND2D1BWP7T $T=101200 357120 0 180 $X=98670 $Y=352910
X1586 79 1 149 201 2 ND2D1BWP7T $T=103440 357120 0 180 $X=100910 $Y=352910
X1587 6 1 226 110 2 ND2D1BWP7T $T=109040 349280 0 0 $X=108750 $Y=349045
X1588 207 1 241 257 2 ND2D1BWP7T $T=137040 357120 0 180 $X=134510 $Y=352910
X1589 1100 1 1065 1098 2 ND2D1BWP7T $T=143760 341440 0 180 $X=141230 $Y=337230
X1590 1099 1 1037 1102 2 ND2D1BWP7T $T=143760 310080 1 0 $X=143470 $Y=305870
X1591 1102 1 992 1108 2 ND2D1BWP7T $T=147120 310080 0 0 $X=146830 $Y=309845
X1592 1098 1 917 1109 2 ND2D1BWP7T $T=168960 333600 1 180 $X=166430 $Y=333365
X1593 335 1 333 332 2 ND2D1BWP7T $T=195280 349280 1 180 $X=192750 $Y=349045
X1594 12 1 20 865 2 872 10 OAI211D1BWP7T $T=23920 333600 0 0 $X=23630 $Y=333365
X1595 1046 1 1048 993 2 1051 917 OAI211D1BWP7T $T=111280 317920 0 0 $X=110990 $Y=317685
X1596 1036 1 1044 1024 2 1053 917 OAI211D1BWP7T $T=111840 325760 0 0 $X=111550 $Y=325525
X1597 1057 1 1062 978 2 243 992 OAI211D1BWP7T $T=129200 302240 0 180 $X=125550 $Y=298030
X1598 1060 1 1023 1055 2 1075 1078 OAI211D1BWP7T $T=128640 325760 1 0 $X=128350 $Y=321550
X1599 405 1 1203 408 2 407 1209 OAI211D1BWP7T $T=258000 294400 0 0 $X=257710 $Y=294165
X1600 1200 1 1204 408 2 1162 1219 OAI211D1BWP7T $T=259120 310080 0 0 $X=258830 $Y=309845
X1601 1210 1 1212 408 2 1164 1213 OAI211D1BWP7T $T=263040 325760 0 0 $X=262750 $Y=325525
X1602 415 1 1214 408 2 1184 1215 OAI211D1BWP7T $T=266400 333600 0 0 $X=266110 $Y=333365
X1603 461 1 1235 1220 2 1237 453 OAI211D1BWP7T $T=294960 349280 0 180 $X=291310 $Y=345070
X1604 1276 1 1277 1278 2 506 437 OAI211D1BWP7T $T=333600 341440 0 0 $X=333310 $Y=341205
X1605 1330 1 1326 1325 2 599 437 OAI211D1BWP7T $T=400800 341440 1 180 $X=397150 $Y=341205
X1606 1340 1 1334 1337 2 1335 437 OAI211D1BWP7T $T=422080 333600 0 180 $X=418430 $Y=329390
X1607 108 2 63 70 18 1 891 NR4D2BWP7T $T=54160 317920 1 180 $X=40990 $Y=317685
X1608 43 2 126 926 1 NR2XD0BWP7T $T=65920 349280 0 0 $X=65630 $Y=349045
X1609 90 2 213 223 1 NR2XD0BWP7T $T=115200 302240 0 180 $X=112670 $Y=298030
X1610 46 1 886 52 12 900 2 ND4D1BWP7T $T=40720 333600 0 0 $X=40430 $Y=333365
X1611 67 1 27 908 60 904 2 ND4D1BWP7T $T=50240 302240 0 180 $X=46030 $Y=298030
X1612 27 1 68 85 88 915 2 ND4D1BWP7T $T=49120 294400 0 0 $X=48830 $Y=294165
X1613 112 1 9 866 117 939 2 ND4D1BWP7T $T=58080 294400 0 0 $X=57790 $Y=294165
X1614 932 1 940 75 866 116 2 ND4D1BWP7T $T=63120 302240 1 180 $X=58910 $Y=302005
X1615 932 1 123 124 54 960 2 ND4D1BWP7T $T=62000 294400 0 0 $X=61710 $Y=294165
X1616 877 1 44 926 143 980 2 ND4D1BWP7T $T=68160 349280 0 0 $X=67870 $Y=349045
X1617 969 1 52 161 155 164 2 ND4D1BWP7T $T=82160 349280 0 0 $X=81870 $Y=349045
X1618 84 1 149 873 162 994 2 ND4D1BWP7T $T=82720 341440 0 0 $X=82430 $Y=341205
X1619 182 1 105 897 189 1019 2 ND4D1BWP7T $T=91120 294400 0 0 $X=90830 $Y=294165
X1620 18 876 923 919 927 1 2 OAI31D1BWP7T $T=51920 325760 1 0 $X=51630 $Y=321550
X1621 234 61 1036 209 911 1 2 OAI31D1BWP7T $T=107360 341440 0 180 $X=103150 $Y=337230
X1622 971 220 1046 233 911 1 2 OAI31D1BWP7T $T=110720 333600 0 0 $X=110430 $Y=333365
X1623 167 236 1057 237 927 1 2 OAI31D1BWP7T $T=121920 302240 1 0 $X=121630 $Y=298030
X1624 235 971 1060 239 212 1 2 OAI31D1BWP7T $T=121920 349280 1 0 $X=121630 $Y=345070
X1625 1016 218 1067 962 248 1 2 OAI31D1BWP7T $T=125840 310080 1 0 $X=125550 $Y=305870
X1626 246 221 1068 1015 212 1 2 OAI31D1BWP7T $T=129760 349280 0 180 $X=125550 $Y=345070
X1627 256 915 1082 1019 240 1 2 OAI31D1BWP7T $T=134240 302240 1 180 $X=130030 $Y=302005
X1628 131 263 1085 894 248 1 2 OAI31D1BWP7T $T=139280 317920 0 180 $X=135070 $Y=313710
X1629 960 266 1093 270 240 1 2 OAI31D1BWP7T $T=139840 302240 1 0 $X=139550 $Y=298030
X1630 268 269 1079 273 226 1 2 OAI31D1BWP7T $T=140960 349280 1 0 $X=140670 $Y=345070
X1631 73 188 869 1006 1004 1 2 AOI31D0BWP7T $T=92240 325760 0 0 $X=91950 $Y=325525
X1632 1030 153 117 1026 1037 1 2 AOI31D0BWP7T $T=103440 310080 1 0 $X=103150 $Y=305870
X1633 228 989 232 1050 975 1 2 AOI31D0BWP7T $T=111280 310080 1 0 $X=110990 $Y=305870
X1634 1061 991 1059 1063 1004 1 2 AOI31D0BWP7T $T=124160 333600 1 0 $X=123870 $Y=329390
X1635 1042 254 143 1081 1065 1 2 AOI31D0BWP7T $T=130880 341440 0 0 $X=130590 $Y=341205
X1636 946 1 122 121 2 942 ND3D0BWP7T $T=64240 349280 1 180 $X=61150 $Y=349045
X1637 136 1 120 944 2 950 ND3D0BWP7T $T=65920 341440 0 180 $X=62830 $Y=337230
X1638 956 1 954 117 2 962 ND3D0BWP7T $T=67040 302240 0 0 $X=66750 $Y=302005
X1639 156 1 149 52 2 938 ND3D0BWP7T $T=82720 341440 1 180 $X=79630 $Y=341205
X1640 29 1 105 202 2 1016 ND3D0BWP7T $T=97840 294400 0 0 $X=97550 $Y=294165
X1641 50 1 2 35 28 888 885 NR4D0BWP7T $T=42400 333600 0 180 $X=38750 $Y=329390
X1642 98 1 2 78 104 905 107 NR4D0BWP7T $T=54160 294400 0 0 $X=53870 $Y=294165
X1643 90 1 2 78 70 956 952 NR4D0BWP7T $T=63120 302240 0 0 $X=62830 $Y=302005
X1644 98 1 2 135 130 954 935 NR4D0BWP7T $T=67600 302240 0 180 $X=63950 $Y=298030
X1645 900 1 2 931 870 964 141 NR4D0BWP7T $T=67040 325760 0 0 $X=66750 $Y=325525
X1646 119 1 2 982 24 986 952 NR4D0BWP7T $T=79920 302240 1 0 $X=79630 $Y=298030
X1647 168 1 2 976 983 984 28 NR4D0BWP7T $T=83280 333600 0 180 $X=79630 $Y=329390
X1648 963 1 2 170 175 998 977 NR4D0BWP7T $T=86640 341440 0 0 $X=86350 $Y=341205
X1649 980 1 2 1013 958 1014 938 NR4D0BWP7T $T=98400 341440 0 180 $X=94750 $Y=337230
X1650 205 1 2 187 199 1012 195 NR4D0BWP7T $T=100080 302240 1 180 $X=96430 $Y=302005
X1651 218 1 2 915 187 1030 196 NR4D0BWP7T $T=104560 302240 0 180 $X=100910 $Y=298030
X1652 219 1 2 221 217 1042 885 NR4D0BWP7T $T=110160 349280 0 180 $X=106510 $Y=345070
X1653 231 1 2 211 173 1043 967 NR4D0BWP7T $T=112960 294400 1 180 $X=109310 $Y=294165
X1654 863 864 2 866 1 NR2D2BWP7T $T=21120 310080 1 0 $X=20830 $Y=305870
X1655 423 421 2 1229 1 NR2D2BWP7T $T=291040 310080 0 0 $X=290750 $Y=309845
X1656 1162 1 2 1159 BUFFD0BWP7T $T=217120 325760 1 180 $X=214590 $Y=325525
X1657 1287 1 2 1285 BUFFD0BWP7T $T=350960 325760 1 180 $X=348430 $Y=325525
X1658 1331 1 2 1325 BUFFD0BWP7T $T=409200 333600 0 180 $X=406670 $Y=329390
X1659 57 943 968 970 975 2 1 AOI31D1BWP7T $T=69280 310080 1 0 $X=68990 $Y=305870
X1660 903 881 988 924 992 2 1 AOI31D1BWP7T $T=82160 317920 0 0 $X=81870 $Y=317685
X1661 998 53 1003 184 1004 2 1 AOI31D1BWP7T $T=90000 341440 0 0 $X=89710 $Y=341205
X1662 1010 891 191 180 975 2 1 AOI31D1BWP7T $T=96160 310080 1 180 $X=91950 $Y=309845
X1663 1043 223 1040 183 1037 2 1 AOI31D1BWP7T $T=111280 310080 0 180 $X=107070 $Y=305870
X1664 1074 1049 1070 242 1065 2 1 AOI31D1BWP7T $T=130320 341440 1 180 $X=126110 $Y=341205
X1665 27 1 9 17 15 867 2 ND4D0BWP7T $T=27840 317920 1 180 $X=24190 $Y=317685
X1666 892 1 888 49 19 896 2 ND4D0BWP7T $T=40720 325760 0 0 $X=40430 $Y=325525
X1667 47 1 893 55 53 901 2 ND4D0BWP7T $T=40720 349280 0 0 $X=40430 $Y=349045
X1668 29 1 898 60 57 879 2 ND4D0BWP7T $T=45760 310080 0 180 $X=42110 $Y=305870
X1669 83 1 80 912 893 907 2 ND4D0BWP7T $T=51360 341440 0 180 $X=47710 $Y=337230
X1670 105 1 102 924 898 919 2 ND4D0BWP7T $T=56960 302240 1 180 $X=53310 $Y=302005
X1671 83 1 103 920 106 930 2 ND4D0BWP7T $T=54160 341440 1 0 $X=53870 $Y=337230
X1672 109 1 120 920 947 937 2 ND4D0BWP7T $T=60880 333600 0 0 $X=60590 $Y=333365
X1673 111 1 129 52 873 963 2 ND4D0BWP7T $T=66480 341440 0 0 $X=66190 $Y=341205
X1674 877 1 136 873 142 966 2 ND4D0BWP7T $T=68160 341440 1 0 $X=67870 $Y=337230
X1675 140 1 940 68 45 979 2 ND4D0BWP7T $T=69840 294400 0 0 $X=69550 $Y=294165
X1676 47 1 969 133 146 976 2 ND4D0BWP7T $T=69840 341440 0 0 $X=69550 $Y=341205
X1677 163 1 124 990 903 987 2 ND4D0BWP7T $T=86640 310080 1 180 $X=82990 $Y=309845
X1678 109 1 83 142 997 1001 2 ND4D0BWP7T $T=86080 341440 1 0 $X=85790 $Y=337230
X1679 109 1 995 174 49 999 2 ND4D0BWP7T $T=86640 325760 0 0 $X=86350 $Y=325525
X1680 922 1 177 178 180 1002 2 ND4D0BWP7T $T=88320 310080 0 0 $X=88030 $Y=309845
X1681 149 1 83 955 1017 1015 2 ND4D0BWP7T $T=95600 341440 0 0 $X=95310 $Y=341205
X1682 918 1 1025 1017 1027 1022 2 ND4D0BWP7T $T=99520 333600 0 0 $X=99230 $Y=333365
X1683 871 1 204 203 1027 1028 2 ND4D0BWP7T $T=99520 349280 1 0 $X=99230 $Y=345070
X1684 1009 1 208 210 1027 1033 2 ND4D0BWP7T $T=102880 349280 1 0 $X=102590 $Y=345070
X1685 224 1 190 902 1020 1031 2 ND4D0BWP7T $T=110160 317920 0 180 $X=106510 $Y=313710
X1686 946 1 225 1041 985 1038 2 ND4D0BWP7T $T=111280 325760 1 180 $X=107630 $Y=325525
X1687 115 1 244 1049 247 1071 2 ND4D0BWP7T $T=127520 349280 0 0 $X=127230 $Y=349045
X1688 965 1 1067 262 1093 1095 2 ND4D0BWP7T $T=136480 310080 1 0 $X=136190 $Y=305870
X1689 48 1 891 2 889 894 IND3D1BWP7T $T=40160 317920 1 0 $X=39870 $Y=313710
X1690 11 864 14 2 1 NR2D1P5BWP7T $T=25040 302240 0 180 $X=20830 $Y=298030
X1691 421 594 595 2 1 NR2D1P5BWP7T $T=399120 317920 1 180 $X=394910 $Y=317685
X1692 866 2 33 876 879 882 1 INR4D0BWP7T $T=26720 325760 1 0 $X=26430 $Y=321550
X1693 111 2 938 872 114 944 1 INR4D0BWP7T $T=57520 341440 1 0 $X=57230 $Y=337230
X1694 210 2 61 220 921 1041 1 INR4D0BWP7T $T=105680 341440 0 0 $X=105390 $Y=341205
X1695 875 1 33 71 903 2 NR3D1BWP7T $T=48000 310080 1 180 $X=43230 $Y=309845
X1696 987 1 151 952 989 2 NR3D1BWP7T $T=80480 317920 1 0 $X=80190 $Y=313710
X1697 125 1 141 157 991 2 NR3D1BWP7T $T=82160 349280 1 0 $X=81870 $Y=345070
X1698 119 1 925 891 951 948 2 IND4D0BWP7T $T=60880 317920 1 0 $X=60590 $Y=313710
X1699 900 1 128 73 941 137 2 IND4D0BWP7T $T=63120 325760 0 0 $X=62830 $Y=325525
X1700 900 1 869 947 973 972 2 IND4D0BWP7T $T=69280 325760 1 0 $X=68990 $Y=321550
X1701 148 1 155 128 1000 984 2 IND4D0BWP7T $T=80480 325760 1 0 $X=80190 $Y=321550
X1702 904 1 1020 925 1029 206 2 IND4D0BWP7T $T=97840 310080 1 0 $X=97550 $Y=305870
X1703 87 1 934 115 931 111 2 IND4D1BWP7T $T=56960 349280 0 0 $X=56670 $Y=349045
X1704 215 874 219 958 2 1 1054 OR4D0BWP7T $T=106800 333600 1 0 $X=106510 $Y=329390
X1705 164 1079 255 169 2 1 1089 OR4D0BWP7T $T=131440 349280 1 0 $X=131150 $Y=345070
X1706 906 86 901 916 926 1 2 INR4D1BWP7T $T=49120 349280 0 0 $X=48830 $Y=349045
X1707 958 983 981 985 47 1 2 INR4D1BWP7T $T=86640 333600 1 180 $X=79630 $Y=333365
X1708 185 93 1007 1009 120 1 2 INR4D1BWP7T $T=91680 357120 1 0 $X=91390 $Y=352910
X1709 14 2 863 1 13 NR2XD1BWP7T $T=28960 302240 0 180 $X=24750 $Y=298030
X1710 865 2 58 1 241 NR2XD1BWP7T $T=121920 357120 1 0 $X=121630 $Y=352910
X1711 1100 2 911 1 1098 NR2XD1BWP7T $T=147680 341440 0 180 $X=143470 $Y=337230
X1712 1102 2 248 1 1108 NR2XD1BWP7T $T=145440 317920 1 0 $X=145150 $Y=313710
X1713 1098 2 1045 1 1109 NR2XD1BWP7T $T=157200 333600 1 180 $X=152990 $Y=333365
X1714 285 2 207 1 296 NR2XD1BWP7T $T=168400 357120 0 180 $X=164190 $Y=352910
X1715 1321 2 611 1 421 NR2XD1BWP7T $T=405280 317920 0 0 $X=404990 $Y=317685
X1716 1077 1 258 259 2 992 1090 OAI211D0BWP7T $T=134240 294400 0 0 $X=133950 $Y=294165
X1717 1086 1 1034 261 2 1078 1097 OAI211D0BWP7T $T=135920 325760 1 0 $X=135630 $Y=321550
X1718 460 1 1239 1186 2 453 1238 OAI211D0BWP7T $T=296640 317920 0 180 $X=292990 $Y=313710
X1719 548 1 1296 1293 2 453 1287 OAI211D0BWP7T $T=358240 325760 0 180 $X=354590 $Y=321550
X1720 12 1 20 10 874 865 2 OAI211D2BWP7T $T=22800 333600 1 0 $X=22510 $Y=329390
X1721 447 1 1228 437 434 1222 2 OAI211D2BWP7T $T=282080 302240 1 180 $X=275630 $Y=302005
X1722 1226 1 1227 437 433 442 2 OAI211D2BWP7T $T=282080 317920 1 180 $X=275630 $Y=317685
X1723 1261 1 1263 482 348 408 2 OAI211D2BWP7T $T=314560 341440 1 180 $X=308110 $Y=341205
X1724 548 1 1302 453 542 1298 2 OAI211D2BWP7T $T=361600 325760 1 180 $X=355150 $Y=325525
X1725 40 99 100 884 1 2 928 AO211D0BWP7T $T=53040 302240 1 0 $X=52750 $Y=298030
X1726 138 2 952 948 99 95 1 AOI211D2BWP7T $T=69280 310080 1 180 $X=62830 $Y=309845
X1727 1070 2 1058 1069 1045 1056 1 AOI211D2BWP7T $T=131440 317920 1 180 $X=124990 $Y=317685
X1728 1099 2 927 1102 1 NR2D3BWP7T $T=142080 310080 0 0 $X=141790 $Y=309845
X1729 268 2 201 278 1 NR2D3BWP7T $T=151040 349280 1 180 $X=145710 $Y=349045
X1730 69 52 4 1 2 ND2D2BWP7T $T=44640 357120 1 0 $X=44350 $Y=352910
X1731 274 273 207 1 2 ND2D2BWP7T $T=155520 349280 1 180 $X=151310 $Y=349045
X1732 950 1 2 870 35 953 NR3D0BWP7T $T=64800 333600 0 0 $X=64510 $Y=333365
X1733 145 1 2 952 967 961 NR3D0BWP7T $T=72080 310080 1 180 $X=68990 $Y=309845
X1734 974 1 2 885 169 995 NR3D0BWP7T $T=86640 333600 0 0 $X=86350 $Y=333365
X1735 193 1 2 171 181 997 NR3D0BWP7T $T=95040 349280 0 180 $X=91950 $Y=345070
X1736 1016 1 2 196 967 194 NR3D0BWP7T $T=98400 302240 0 180 $X=95310 $Y=298030
X1737 198 1022 1 1006 1023 2 AOI21D1BWP7T $T=102320 325760 0 180 $X=98670 $Y=321550
X1738 535 1286 1 1290 1279 2 AOI21D1BWP7T $T=349280 333600 1 0 $X=348990 $Y=329390
X1739 880 873 886 47 64 1 2 ND4D2BWP7T $T=39040 341440 1 0 $X=38750 $Y=337230
X1740 77 5 75 889 90 1 2 ND4D2BWP7T $T=53040 310080 0 180 $X=45470 $Y=305870
X1741 899 92 886 81 921 1 2 ND4D2BWP7T $T=50240 341440 0 0 $X=49950 $Y=341205
X1742 961 127 66 932 131 1 2 ND4D2BWP7T $T=67040 317920 1 180 $X=59470 $Y=317685
X1743 926 92 129 134 949 1 2 ND4D2BWP7T $T=60320 357120 1 0 $X=60030 $Y=352910
X1744 155 916 122 192 1005 1 2 ND4D2BWP7T $T=88320 349280 0 0 $X=88030 $Y=349045
X1745 1091 1076 275 1096 272 1 2 ND4D2BWP7T $T=139840 333600 1 0 $X=139550 $Y=329390
X1746 927 1 965 951 139 98 2 OAI31D2BWP7T $T=72080 317920 0 180 $X=65070 $Y=313710
X1747 198 1 1008 999 193 168 2 OAI31D2BWP7T $T=97280 325760 0 180 $X=90270 $Y=321550
X1748 1045 1 1076 909 251 959 2 OAI31D2BWP7T $T=133120 325760 1 180 $X=126110 $Y=325525
X1749 247 1 1066 865 264 274 2 OAI31D2BWP7T $T=137040 357120 1 0 $X=136750 $Y=352910
X1750 1045 1 1106 996 974 219 2 OAI31D2BWP7T $T=152160 333600 1 180 $X=145150 $Y=333365
X1751 38 1 52 59 2 61 ND3D1BWP7T $T=40720 357120 1 0 $X=40430 $Y=352910
X1752 31 1 68 905 2 72 ND3D1BWP7T $T=44640 294400 0 0 $X=44350 $Y=294165
X1753 109 1 132 953 2 959 ND3D1BWP7T $T=64240 333600 1 0 $X=63950 $Y=329390
X1754 47 1 83 103 2 974 ND3D1BWP7T $T=69840 333600 0 0 $X=69550 $Y=333365
X1755 147 1 165 166 2 996 ND3D1BWP7T $T=84400 357120 1 0 $X=84110 $Y=352910
X1756 264 1 110 257 2 946 ND3D1BWP7T $T=139280 349280 1 180 $X=135630 $Y=349045
X1757 72 2 70 91 1 908 95 AOI211D1BWP7T $T=50240 302240 0 0 $X=49950 $Y=302005
X1758 107 2 935 113 1 943 95 AOI211D1BWP7T $T=58640 310080 1 0 $X=58350 $Y=305870
X1759 1244 2 1245 464 1 1239 395 AOI211D1BWP7T $T=300000 317920 0 180 $X=296350 $Y=313710
X1760 1274 2 1229 510 1 1273 397 AOI211D1BWP7T $T=333600 325760 0 0 $X=333310 $Y=325525
X1761 613 2 594 614 1 1334 397 AOI211D1BWP7T $T=415920 317920 0 0 $X=415630 $Y=317685
X1762 629 2 611 1344 1 1343 397 AOI211D1BWP7T $T=426000 325760 0 180 $X=422350 $Y=321550
X1763 94 1 172 163 982 140 2 IND4D2BWP7T $T=92240 302240 0 180 $X=83550 $Y=298030
X1764 133 2 920 125 1 INR2D1BWP7T $T=66480 341440 1 180 $X=63390 $Y=341205
X1793 1 2 ICV_19 $T=27840 317920 0 0 $X=27550 $Y=317685
X1794 1 2 ICV_19 $T=35120 325760 1 0 $X=34830 $Y=321550
X1795 1 2 ICV_19 $T=144880 349280 1 0 $X=144590 $Y=345070
X1796 1 2 ICV_19 $T=146000 341440 0 0 $X=145710 $Y=341205
X1797 1 2 ICV_19 $T=178480 341440 1 0 $X=178190 $Y=337230
X1798 1 2 ICV_19 $T=179600 325760 0 0 $X=179310 $Y=325525
X1799 1 2 ICV_19 $T=195840 302240 1 0 $X=195550 $Y=298030
X1800 1 2 ICV_19 $T=222160 349280 1 0 $X=221870 $Y=345070
X1801 1 2 ICV_19 $T=237840 349280 0 0 $X=237550 $Y=349045
X1802 1 2 ICV_19 $T=264160 341440 1 0 $X=263870 $Y=337230
X1803 1 2 ICV_19 $T=279840 349280 0 0 $X=279550 $Y=349045
X1804 1 2 ICV_19 $T=309520 341440 1 0 $X=309230 $Y=337230
X1805 1 2 ICV_19 $T=313440 333600 0 0 $X=313150 $Y=333365
X1806 1 2 ICV_19 $T=321840 333600 1 0 $X=321550 $Y=329390
X1807 1 2 ICV_19 $T=321840 349280 1 0 $X=321550 $Y=345070
X1808 1 2 ICV_19 $T=378960 317920 0 0 $X=378670 $Y=317685
X1809 1 2 ICV_19 $T=380080 349280 0 0 $X=379790 $Y=349045
X1810 1 2 ICV_19 $T=398560 310080 0 0 $X=398270 $Y=309845
X1811 1 2 ICV_19 $T=437760 333600 1 0 $X=437470 $Y=329390
X1812 1 2 ICV_19 $T=447840 349280 1 0 $X=447550 $Y=345070
X1813 1 2 ICV_21 $T=152720 341440 1 0 $X=152430 $Y=337230
X1814 1 2 ICV_21 $T=219920 294400 0 0 $X=219630 $Y=294165
X1815 1 2 ICV_21 $T=255760 310080 1 0 $X=255470 $Y=305870
X1816 1 2 ICV_21 $T=266400 325760 0 0 $X=266110 $Y=325525
X1817 1 2 ICV_21 $T=278720 333600 0 0 $X=278430 $Y=333365
X1818 1 2 ICV_21 $T=320720 341440 1 0 $X=320430 $Y=337230
X1819 1 2 ICV_21 $T=338080 310080 0 0 $X=337790 $Y=309845
X1820 1 2 ICV_21 $T=346480 341440 0 0 $X=346190 $Y=341205
X1821 1 2 ICV_21 $T=362720 317920 1 0 $X=362430 $Y=313710
X1822 1 2 ICV_21 $T=362720 317920 0 0 $X=362430 $Y=317685
X1823 1 2 ICV_21 $T=382880 333600 1 0 $X=382590 $Y=329390
X1824 1 2 ICV_21 $T=391280 349280 0 0 $X=390990 $Y=349045
X1825 1 2 ICV_21 $T=404720 302240 1 0 $X=404430 $Y=298030
X1826 1 2 ICV_21 $T=404720 302240 0 0 $X=404430 $Y=302005
X1827 1 2 ICV_21 $T=404720 357120 1 0 $X=404430 $Y=352910
X1828 1 2 ICV_21 $T=413120 310080 0 0 $X=412830 $Y=309845
X1829 1 2 ICV_21 $T=424880 341440 1 0 $X=424590 $Y=337230
X1830 1 2 ICV_21 $T=432720 325760 1 0 $X=432430 $Y=321550
X1831 1 2 ICV_21 $T=434400 333600 0 0 $X=434110 $Y=333365
X1832 1 2 ICV_21 $T=434960 341440 1 0 $X=434670 $Y=337230
X1837 314 1180 303 1365 2 1 365 DFCND1BWP7T $T=237280 310080 1 180 $X=224110 $Y=309845
X1838 314 372 303 1366 2 1 389 DFCND1BWP7T $T=227200 294400 0 0 $X=226910 $Y=294165
X1839 314 1177 303 1367 2 1 369 DFCND1BWP7T $T=240080 310080 0 180 $X=226910 $Y=305870
X1840 314 1190 303 1368 2 1 1195 DFCND1BWP7T $T=248480 317920 0 0 $X=248190 $Y=317685
X1841 314 1194 303 1369 2 1 1193 DFCND1BWP7T $T=249600 349280 1 0 $X=249310 $Y=345070
X1842 314 1198 403 1370 2 1 368 DFCND1BWP7T $T=263040 357120 0 180 $X=249870 $Y=352910
X1843 314 1189 403 1371 2 1 1192 DFCND1BWP7T $T=264160 341440 0 180 $X=250990 $Y=337230
X1844 314 404 403 414 2 1 416 DFCND1BWP7T $T=254640 302240 1 0 $X=254350 $Y=298030
X1845 530 1284 523 1292 2 1 1297 DFCND1BWP7T $T=345360 310080 0 0 $X=345070 $Y=309845
X1846 530 1295 523 1372 2 1 1205 DFCND1BWP7T $T=359360 349280 0 180 $X=346190 $Y=345070
X1847 910 1 2 35 110 1018 207 AOI211XD0BWP7T $T=98960 349280 0 0 $X=98670 $Y=349045
X1848 1040 1 2 1064 1002 1072 248 AOI211XD0BWP7T $T=127520 317920 1 0 $X=127230 $Y=313710
X1849 1230 1 2 1229 448 1227 397 AOI211XD0BWP7T $T=282640 310080 1 180 $X=278990 $Y=309845
X1850 1236 1 2 1234 455 1228 397 AOI211XD0BWP7T $T=294960 302240 1 180 $X=291310 $Y=302005
X1851 1258 1 2 1234 1249 1252 397 AOI211XD0BWP7T $T=306720 302240 1 180 $X=303070 $Y=302005
X1852 1279 1 2 1229 507 1277 397 AOI211XD0BWP7T $T=336960 333600 1 180 $X=333310 $Y=333365
X1853 1312 1 2 1310 1309 1308 395 AOI211XD0BWP7T $T=377840 333600 0 180 $X=374190 $Y=329390
X1854 1342 1 2 611 1332 1326 397 AOI211XD0BWP7T $T=422640 341440 1 180 $X=418990 $Y=341205
X1855 314 1211 403 1373 409 1 2 DFCND2BWP7T $T=261360 325760 1 0 $X=261070 $Y=321550
X1856 530 1306 523 584 1301 1 2 DFCND2BWP7T $T=377280 349280 1 0 $X=376990 $Y=345070
X1857 871 1 22 865 10 2 OAI21D2BWP7T $T=27840 349280 0 180 $X=22510 $Y=345070
X1858 1225 1 1150 439 1223 2 OAI21D2BWP7T $T=280400 349280 0 180 $X=275070 $Y=345070
X1859 1240 1 1166 439 456 2 OAI21D2BWP7T $T=296640 341440 0 180 $X=291310 $Y=337230
X1860 1248 1 1165 439 1243 2 OAI21D2BWP7T $T=302240 333600 0 180 $X=296910 $Y=329390
X1861 1262 1 1153 439 1260 2 OAI21D2BWP7T $T=313440 333600 1 180 $X=308110 $Y=333365
X1862 1269 1 1132 439 1266 2 OAI21D2BWP7T $T=320720 341440 0 180 $X=315390 $Y=337230
X1863 498 1 1135 439 1268 2 OAI21D2BWP7T $T=321840 333600 0 180 $X=316510 $Y=329390
X1864 1316 1 1144 551 1315 2 OAI21D2BWP7T $T=380080 349280 1 180 $X=374750 $Y=349045
X1865 1289 361 1 1137 531 2 IOA21D1BWP7T $T=349840 317920 1 180 $X=346190 $Y=317685
X1866 478 437 1 474 2 1258 1254 OAI22D1BWP7T $T=308960 294400 1 180 $X=304750 $Y=294165
X1867 1187 437 1 474 2 1251 1257 OAI22D1BWP7T $T=310080 310080 1 180 $X=305870 $Y=309845
X1868 1267 437 1 474 2 1274 1264 OAI22D1BWP7T $T=321280 310080 0 0 $X=320990 $Y=309845
X1869 1300 474 1 437 2 558 1304 OAI22D1BWP7T $T=363280 341440 0 0 $X=362990 $Y=341205
X1870 1322 437 1 474 2 598 1329 OAI22D1BWP7T $T=400800 357120 1 0 $X=400510 $Y=352910
X1871 668 1 2 706 DEL1BWP7T $T=465200 317920 1 0 $X=464910 $Y=313710
X1872 1148 576 1356 1197 683 1 2 687 AO221D1BWP7T $T=461280 317920 0 0 $X=460990 $Y=317685
X1873 314 1161 303 1374 2 1 1168 DFCND0BWP7T $T=210960 333600 1 0 $X=210670 $Y=329390
X1874 314 1179 303 1375 2 1 1172 DFCND0BWP7T $T=233920 341440 0 180 $X=220750 $Y=337230
X1875 314 1176 303 1376 2 1 1182 DFCND0BWP7T $T=222720 349280 0 0 $X=222430 $Y=349045
X1876 314 1171 303 1377 2 1 1175 DFCND0BWP7T $T=236160 325760 0 180 $X=222990 $Y=321550
X1877 314 379 303 1378 2 1 1170 DFCND0BWP7T $T=238400 302240 0 180 $X=225230 $Y=298030
X1878 314 1183 303 1379 2 1 1178 DFCND0BWP7T $T=239520 333600 1 180 $X=226350 $Y=333365
X1879 314 1191 303 1208 2 1 401 DFCND0BWP7T $T=249040 325760 0 0 $X=248750 $Y=325525
X1880 544 541 523 1380 2 1 512 DFCND0BWP7T $T=358240 357120 0 180 $X=345070 $Y=352910
X1881 530 1288 523 1299 2 1 1303 DFCND0BWP7T $T=348720 310080 1 0 $X=348430 $Y=305870
X1882 530 1320 523 1324 2 1 1294 DFCND0BWP7T $T=382320 341440 0 0 $X=382030 $Y=341205
X1883 530 592 523 604 2 1 1328 DFCND0BWP7T $T=392400 294400 0 0 $X=392110 $Y=294165
X1884 530 632 523 1338 2 1 1339 DFCND0BWP7T $T=433840 294400 1 180 $X=420670 $Y=294165
X1885 553 551 418 549 538 1292 2 1291 1 OA222D0BWP7T $T=362160 302240 1 180 $X=355710 $Y=302005
X1886 610 551 418 606 538 1324 2 1323 1 OA222D0BWP7T $T=406400 333600 1 180 $X=399950 $Y=333365
X1887 628 551 418 621 538 620 2 1336 1 OA222D0BWP7T $T=425440 349280 1 180 $X=418990 $Y=349045
X1888 1021 2 968 1 1032 927 1031 AOI211XD1BWP7T $T=97840 317920 1 0 $X=97550 $Y=313710
X1889 1088 2 1073 1 1101 911 1005 AOI211XD1BWP7T $T=135360 333600 0 0 $X=135070 $Y=333365
X1890 528 555 1 2 INVD2P5BWP7T $T=381200 317920 0 180 $X=378110 $Y=313710
X1891 474 398 1 2 INVD6BWP7T $T=308960 317920 0 180 $X=303630 $Y=313710
X1892 524 551 1 2 INVD6BWP7T $T=435520 357120 1 0 $X=435230 $Y=352910
X1893 551 555 1 418 543 538 1292 2 1288 OAI222D2BWP7T $T=362720 317920 0 180 $X=352350 $Y=313710
X1894 551 634 1 418 621 538 626 2 624 OAI222D2BWP7T $T=432720 349280 0 180 $X=422350 $Y=345070
X1895 1238 451 450 1 2 XOR2D2BWP7T $T=296640 317920 1 180 $X=289630 $Y=317685
X1896 245 72 250 1077 927 1 2 OAI31D0BWP7T $T=129200 294400 0 0 $X=128910 $Y=294165
X1897 367 418 1 2 CKND4BWP7T $T=270880 349280 1 180 $X=266670 $Y=349045
X1898 36 29 40 1 2 ND2D1P5BWP7T $T=30640 294400 1 180 $X=26430 $Y=294165
X1899 279 278 269 1 2 ND2D1P5BWP7T $T=151600 333600 1 0 $X=151310 $Y=329390
X1900 107 88 925 929 1 2 63 IIND4D1BWP7T $T=58640 310080 1 180 $X=52750 $Y=309845
X1901 683 665 1 2 CKND6BWP7T $T=467440 325760 1 180 $X=462110 $Y=325525
X1902 665 1 672 402 1360 685 2 681 OAI221D2BWP7T $T=459040 357120 1 0 $X=458750 $Y=352910
X1903 665 1 487 326 692 1361 2 1362 OAI221D2BWP7T $T=469680 302240 1 180 $X=460430 $Y=302005
X1904 1 2 ICV_23 $T=119120 310080 1 0 $X=118830 $Y=305870
X1905 1 2 ICV_23 $T=153280 349280 1 0 $X=152990 $Y=345070
X1906 1 2 ICV_23 $T=153280 357120 1 0 $X=152990 $Y=352910
X1907 1 2 ICV_23 $T=161120 349280 0 0 $X=160830 $Y=349045
X1908 1 2 ICV_23 $T=181840 310080 0 0 $X=181550 $Y=309845
X1909 1 2 ICV_23 $T=195280 317920 0 0 $X=194990 $Y=317685
X1910 1 2 ICV_23 $T=195280 341440 0 0 $X=194990 $Y=341205
X1911 1 2 ICV_23 $T=195280 349280 0 0 $X=194990 $Y=349045
X1912 1 2 ICV_23 $T=237280 310080 0 0 $X=236990 $Y=309845
X1913 1 2 ICV_23 $T=294960 302240 0 0 $X=294670 $Y=302005
X1914 1 2 ICV_23 $T=296640 317920 0 0 $X=296350 $Y=317685
X1915 1 2 ICV_23 $T=329120 325760 1 0 $X=328830 $Y=321550
X1916 1 2 ICV_23 $T=338080 349280 1 0 $X=337790 $Y=345070
X1917 1 2 ICV_23 $T=353760 341440 1 0 $X=353470 $Y=337230
X1918 1 2 ICV_23 $T=361600 294400 0 0 $X=361310 $Y=294165
X1919 1 2 ICV_23 $T=361600 333600 1 0 $X=361310 $Y=329390
X1920 1 2 ICV_23 $T=371120 302240 1 0 $X=370830 $Y=298030
X1921 1 2 ICV_23 $T=371120 310080 1 0 $X=370830 $Y=305870
X1922 1 2 ICV_23 $T=403600 325760 1 0 $X=403310 $Y=321550
X1923 1 2 ICV_23 $T=403600 349280 0 0 $X=403310 $Y=349045
X1924 1 2 ICV_23 $T=405280 294400 0 0 $X=404990 $Y=294165
X1925 1 2 ICV_23 $T=413120 302240 1 0 $X=412830 $Y=298030
X1926 1 2 ICV_23 $T=422080 302240 1 0 $X=421790 $Y=298030
X1927 1 2 ICV_23 $T=433840 341440 0 0 $X=433550 $Y=341205
X1928 1 2 ICV_23 $T=447280 302240 0 0 $X=446990 $Y=302005
X1929 1 2 ICV_23 $T=447280 317920 0 0 $X=446990 $Y=317685
X1930 426 408 1 2 INVD8BWP7T $T=273680 325760 0 0 $X=273390 $Y=325525
X1931 339 530 1 2 INVD8BWP7T $T=354880 294400 0 0 $X=354590 $Y=294165
X1932 289 282 277 297 1 2 1120 AO22D0BWP7T $T=163920 294400 0 0 $X=163630 $Y=294165
X1933 501 487 469 481 1 2 1253 AO22D0BWP7T $T=320720 317920 0 180 $X=315950 $Y=313710
X1934 465 2 469 1 CKND10BWP7T $T=298320 349280 0 0 $X=298030 $Y=349045
X1935 296 257 285 2 304 1 ND3D3BWP7T $T=172320 349280 1 0 $X=172030 $Y=345070
X1936 1122 257 296 79 1 2 AN3D2BWP7T $T=168960 349280 0 180 $X=164190 $Y=345070
X1937 269 279 268 865 2 1 OR3D2BWP7T $T=148240 357120 0 180 $X=143470 $Y=352910
X1938 1084 1069 1025 1087 1078 1069 2 1 AOI32D1BWP7T $T=135920 317920 1 180 $X=131150 $Y=317685
X1939 1035 1101 991 1104 917 1101 2 1 AOI32D1BWP7T $T=148240 325760 1 180 $X=143470 $Y=325525
X1940 878 45 5 29 2 42 1 ND4D3BWP7T $T=36800 302240 0 0 $X=36510 $Y=302005
X1941 1080 1103 1106 1094 2 276 1 ND4D3BWP7T $T=142640 317920 0 0 $X=142350 $Y=317685
X1942 62 1 73 899 909 2 IND3D2BWP7T $T=44080 325760 0 0 $X=43790 $Y=325525
X1943 16 1 26 873 2 CKND2D2BWP7T $T=25040 349280 0 0 $X=24750 $Y=349045
.ENDS
***************************************
.SUBCKT ICV_25
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT AO221D2BWP7T A2 A1 B2 B1 C Z VSS VDD
** N=13 EP=8 IP=0 FDC=14
M0 12 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=660 $Y=345 $D=0
M1 11 A1 12 VSS N L=1.8e-07 W=1e-06 $X=1260 $Y=345 $D=0
M2 13 B2 VSS VSS N L=1.8e-07 W=1e-06 $X=2910 $Y=345 $D=0
M3 11 B1 13 VSS N L=1.8e-07 W=1e-06 $X=3630 $Y=345 $D=0
M4 VSS C 11 VSS N L=1.8e-07 W=1e-06 $X=4350 $Y=345 $D=0
M5 Z 11 VSS VSS N L=1.8e-07 W=1e-06 $X=5200 $Y=345 $D=0
M6 VSS 11 Z VSS N L=1.8e-07 W=1e-06 $X=5920 $Y=345 $D=0
M7 11 A2 9 VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M8 9 A1 11 VDD P L=1.8e-07 W=1.37e-06 $X=1380 $Y=2205 $D=16
M9 9 B2 10 VDD P L=1.8e-07 W=1.37e-06 $X=2910 $Y=2205 $D=16
M10 10 B1 9 VDD P L=1.8e-07 W=1.37e-06 $X=3630 $Y=2205 $D=16
M11 VDD C 10 VDD P L=1.8e-07 W=1.37e-06 $X=4350 $Y=2205 $D=16
M12 Z 11 VDD VDD P L=1.8e-07 W=1.37e-06 $X=5200 $Y=2205 $D=16
M13 VDD 11 Z VDD P L=1.8e-07 W=1.37e-06 $X=5920 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_26 1 2
** N=2 EP=2 IP=4 FDC=10
X0 1 2 DCAP8BWP7T $T=0 0 0 0 $X=-290 $Y=-235
X1 1 2 ICV_13 $T=4480 0 0 0 $X=4190 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_27 1 2
** N=2 EP=2 IP=4 FDC=4
X1 1 2 ICV_13 $T=1120 0 0 0 $X=830 $Y=-235
.ENDS
***************************************
.SUBCKT OAI22D2BWP7T B1 VSS B2 ZN A1 A2 VDD
** N=12 EP=7 IP=0 FDC=16
M0 VSS B2 8 VSS N L=1.8e-07 W=1e-06 $X=630 $Y=345 $D=0
M1 8 B1 VSS VSS N L=1.8e-07 W=1e-06 $X=1400 $Y=345 $D=0
M2 VSS B1 8 VSS N L=1.8e-07 W=1e-06 $X=2120 $Y=345 $D=0
M3 8 B2 VSS VSS N L=1.8e-07 W=1e-06 $X=2920 $Y=345 $D=0
M4 ZN A2 8 VSS N L=1.8e-07 W=1e-06 $X=3680 $Y=345 $D=0
M5 8 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=4420 $Y=345 $D=0
M6 ZN A1 8 VSS N L=1.8e-07 W=1e-06 $X=5140 $Y=345 $D=0
M7 8 A2 ZN VSS N L=1.8e-07 W=1e-06 $X=5860 $Y=345 $D=0
M8 9 B2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=630 $Y=2205 $D=16
M9 ZN B1 9 VDD P L=1.8e-07 W=1.37e-06 $X=1400 $Y=2205 $D=16
M10 10 B1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2120 $Y=2205 $D=16
M11 VDD B2 10 VDD P L=1.8e-07 W=1.37e-06 $X=2760 $Y=2205 $D=16
M12 11 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3720 $Y=2205 $D=16
M13 ZN A1 11 VDD P L=1.8e-07 W=1.37e-06 $X=4320 $Y=2205 $D=16
M14 12 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=5080 $Y=2205 $D=16
M15 VDD A2 12 VDD P L=1.8e-07 W=1.37e-06 $X=5680 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OAI22D0BWP7T B2 A1 ZN A2 B1 VDD VSS
** N=10 EP=7 IP=0 FDC=8
M0 8 B2 VSS VSS N L=1.8e-07 W=5e-07 $X=625 $Y=480 $D=0
M1 ZN A1 8 VSS N L=1.8e-07 W=5e-07 $X=1225 $Y=735 $D=0
M2 8 A2 ZN VSS N L=1.8e-07 W=5e-07 $X=1945 $Y=735 $D=0
M3 VSS B1 8 VSS N L=1.8e-07 W=5e-07 $X=2555 $Y=345 $D=0
M4 9 B2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=625 $Y=2890 $D=16
M5 ZN B1 9 VDD P L=1.8e-07 W=6.85e-07 $X=1330 $Y=2890 $D=16
M6 10 A1 ZN VDD P L=1.8e-07 W=6.85e-07 $X=2130 $Y=2890 $D=16
M7 VDD A2 10 VDD P L=1.8e-07 W=6.85e-07 $X=2560 $Y=2890 $D=16
.ENDS
***************************************
.SUBCKT BUFFD4BWP7T I Z VSS VDD
** N=5 EP=4 IP=0 FDC=12
M0 5 I VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS I 5 VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=2080 $Y=345 $D=0
M3 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=2800 $Y=345 $D=0
M4 Z 5 VSS VSS N L=1.8e-07 W=1e-06 $X=3520 $Y=345 $D=0
M5 VSS 5 Z VSS N L=1.8e-07 W=1e-06 $X=4240 $Y=345 $D=0
M6 5 I VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M7 VDD I 5 VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M8 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2080 $Y=2205 $D=16
M9 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=2800 $Y=2205 $D=16
M10 Z 5 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3520 $Y=2205 $D=16
M11 VDD 5 Z VDD P L=1.8e-07 W=1.37e-06 $X=4240 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR3D3BWP7T A3 VDD A2 A1 VSS ZN
** N=8 EP=6 IP=0 FDC=30
M0 ZN A3 VSS VSS N L=1.8e-07 W=6e-07 $X=780 $Y=345 $D=0
M1 VSS A3 ZN VSS N L=1.8e-07 W=6e-07 $X=1500 $Y=345 $D=0
M2 ZN A3 VSS VSS N L=1.8e-07 W=6e-07 $X=2220 $Y=345 $D=0
M3 VSS A3 ZN VSS N L=1.8e-07 W=6e-07 $X=2940 $Y=345 $D=0
M4 ZN A3 VSS VSS N L=1.8e-07 W=6e-07 $X=3660 $Y=345 $D=0
M5 VSS A2 ZN VSS N L=1.8e-07 W=6e-07 $X=4380 $Y=345 $D=0
M6 ZN A2 VSS VSS N L=1.8e-07 W=6e-07 $X=5100 $Y=345 $D=0
M7 VSS A2 ZN VSS N L=1.8e-07 W=6e-07 $X=5820 $Y=345 $D=0
M8 ZN A2 VSS VSS N L=1.8e-07 W=6e-07 $X=6540 $Y=345 $D=0
M9 VSS A2 ZN VSS N L=1.8e-07 W=6e-07 $X=7260 $Y=345 $D=0
M10 ZN A1 VSS VSS N L=1.8e-07 W=6e-07 $X=7980 $Y=345 $D=0
M11 VSS A1 ZN VSS N L=1.8e-07 W=6e-07 $X=8700 $Y=345 $D=0
M12 ZN A1 VSS VSS N L=1.8e-07 W=6e-07 $X=9420 $Y=345 $D=0
M13 VSS A1 ZN VSS N L=1.8e-07 W=6e-07 $X=10140 $Y=345 $D=0
M14 ZN A1 VSS VSS N L=1.8e-07 W=6e-07 $X=10860 $Y=345 $D=0
M15 7 A3 VDD VDD P L=1.8e-07 W=1.36e-06 $X=780 $Y=2215 $D=16
M16 VDD A3 7 VDD P L=1.8e-07 W=1.715e-06 $X=1500 $Y=1860 $D=16
M17 7 A3 VDD VDD P L=1.8e-07 W=1.715e-06 $X=2220 $Y=1860 $D=16
M18 VDD A3 7 VDD P L=1.8e-07 W=1.715e-06 $X=2940 $Y=1860 $D=16
M19 7 A3 VDD VDD P L=1.8e-07 W=1.715e-06 $X=3660 $Y=1860 $D=16
M20 8 A2 7 VDD P L=1.8e-07 W=1.645e-06 $X=4380 $Y=1930 $D=16
M21 7 A2 8 VDD P L=1.8e-07 W=1.645e-06 $X=5100 $Y=1930 $D=16
M22 8 A2 7 VDD P L=1.8e-07 W=1.645e-06 $X=5820 $Y=1930 $D=16
M23 7 A2 8 VDD P L=1.8e-07 W=1.645e-06 $X=6540 $Y=1930 $D=16
M24 8 A2 7 VDD P L=1.8e-07 W=1.645e-06 $X=7260 $Y=1930 $D=16
M25 ZN A1 8 VDD P L=1.8e-07 W=1.715e-06 $X=7980 $Y=1860 $D=16
M26 8 A1 ZN VDD P L=1.8e-07 W=1.715e-06 $X=8700 $Y=1860 $D=16
M27 ZN A1 8 VDD P L=1.8e-07 W=1.715e-06 $X=9420 $Y=1860 $D=16
M28 8 A1 ZN VDD P L=1.8e-07 W=1.715e-06 $X=10140 $Y=1860 $D=16
M29 ZN A1 8 VDD P L=1.8e-07 W=1.36e-06 $X=10860 $Y=2215 $D=16
.ENDS
***************************************
.SUBCKT ND4D4BWP7T A1 A2 A3 ZN VSS A4 VDD
** N=10 EP=7 IP=0 FDC=32
M0 ZN A1 8 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 8 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 ZN A1 8 VSS N L=1.8e-07 W=1e-06 $X=2060 $Y=345 $D=0
M3 8 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=2780 $Y=345 $D=0
M4 9 A2 8 VSS N L=1.8e-07 W=1e-06 $X=3500 $Y=345 $D=0
M5 8 A2 9 VSS N L=1.8e-07 W=1e-06 $X=4220 $Y=345 $D=0
M6 9 A2 8 VSS N L=1.8e-07 W=1e-06 $X=4940 $Y=345 $D=0
M7 8 A2 9 VSS N L=1.8e-07 W=1e-06 $X=5660 $Y=345 $D=0
M8 9 A3 10 VSS N L=1.8e-07 W=1e-06 $X=7040 $Y=345 $D=0
M9 10 A3 9 VSS N L=1.8e-07 W=1e-06 $X=7760 $Y=345 $D=0
M10 9 A3 10 VSS N L=1.8e-07 W=1e-06 $X=8480 $Y=345 $D=0
M11 10 A3 9 VSS N L=1.8e-07 W=1e-06 $X=9200 $Y=345 $D=0
M12 VSS A4 10 VSS N L=1.8e-07 W=1e-06 $X=9920 $Y=345 $D=0
M13 10 A4 VSS VSS N L=1.8e-07 W=1e-06 $X=10640 $Y=345 $D=0
M14 VSS A4 10 VSS N L=1.8e-07 W=1e-06 $X=11360 $Y=345 $D=0
M15 10 A4 VSS VSS N L=1.8e-07 W=1e-06 $X=12080 $Y=345 $D=0
M16 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M17 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M18 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M19 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M20 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3500 $Y=2205 $D=16
M21 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4220 $Y=2205 $D=16
M22 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4940 $Y=2205 $D=16
M23 VDD A2 ZN VDD P L=1.8e-07 W=1.36e-06 $X=5660 $Y=2215 $D=16
M24 ZN A3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=7040 $Y=2205 $D=16
M25 VDD A3 ZN VDD P L=1.8e-07 W=1.37e-06 $X=7760 $Y=2205 $D=16
M26 ZN A3 VDD VDD P L=1.8e-07 W=1.37e-06 $X=8480 $Y=2205 $D=16
M27 VDD A3 ZN VDD P L=1.8e-07 W=1.37e-06 $X=9200 $Y=2205 $D=16
M28 ZN A4 VDD VDD P L=1.8e-07 W=1.37e-06 $X=9920 $Y=2205 $D=16
M29 VDD A4 ZN VDD P L=1.8e-07 W=1.37e-06 $X=10640 $Y=2205 $D=16
M30 ZN A4 VDD VDD P L=1.8e-07 W=1.37e-06 $X=11360 $Y=2205 $D=16
M31 VDD A4 ZN VDD P L=1.8e-07 W=1.37e-06 $X=12080 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IOA22D2BWP7T A1 A2 ZN B2 VDD B1 VSS
** N=12 EP=7 IP=0 FDC=14
M0 9 10 VSS VSS N L=1.8e-07 W=1e-06 $X=660 $Y=345 $D=0
M1 11 A1 9 VSS N L=1.8e-07 W=1e-06 $X=1595 $Y=345 $D=0
M2 VSS A2 11 VSS N L=1.8e-07 W=1e-06 $X=2140 $Y=345 $D=0
M3 ZN 9 VSS VSS N L=1.8e-07 W=1e-06 $X=3235 $Y=345 $D=0
M4 VSS 9 ZN VSS N L=1.8e-07 W=1e-06 $X=3955 $Y=345 $D=0
M5 10 B2 VSS VSS N L=1.8e-07 W=5e-07 $X=4640 $Y=845 $D=0
M6 VSS B1 10 VSS N L=1.8e-07 W=5e-07 $X=5360 $Y=845 $D=0
M7 8 10 9 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M8 VDD A1 8 VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M9 8 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2070 $Y=2205 $D=16
M10 ZN 9 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3345 $Y=2205 $D=16
M11 VDD 9 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4065 $Y=2205 $D=16
M12 12 B2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=4805 $Y=2205 $D=16
M13 10 B1 12 VDD P L=1.8e-07 W=1.37e-06 $X=5360 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT CKND8BWP7T I ZN VSS VDD
** N=4 EP=4 IP=0 FDC=15
M0 ZN I VSS VSS N L=1.8e-07 W=7e-07 $X=2080 $Y=345 $D=0
M1 VSS I ZN VSS N L=1.8e-07 W=7e-07 $X=2800 $Y=345 $D=0
M2 ZN I VSS VSS N L=1.8e-07 W=7e-07 $X=3520 $Y=345 $D=0
M3 VSS I ZN VSS N L=1.8e-07 W=7e-07 $X=4240 $Y=345 $D=0
M4 ZN I VSS VSS N L=1.8e-07 W=7e-07 $X=4960 $Y=345 $D=0
M5 VSS I ZN VSS N L=1.8e-07 W=7e-07 $X=5680 $Y=345 $D=0
M6 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=640 $Y=2205 $D=16
M7 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=1360 $Y=2205 $D=16
M8 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=2080 $Y=2205 $D=16
M9 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=2800 $Y=2205 $D=16
M10 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=3520 $Y=2205 $D=16
M11 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=4240 $Y=2205 $D=16
M12 ZN I VDD VDD P L=1.8e-07 W=1.37e-06 $X=4960 $Y=2205 $D=16
M13 VDD I ZN VDD P L=1.8e-07 W=1.37e-06 $X=5680 $Y=2205 $D=16
D14 VSS I DN AREA=2.037e-13 PJ=1.81e-06 $X=140 $Y=860 $D=32
.ENDS
***************************************
.SUBCKT AN2D2BWP7T A1 A2 Z VSS VDD
** N=7 EP=5 IP=0 FDC=8
M0 7 A1 6 VSS N L=1.8e-07 W=1e-06 $X=740 $Y=345 $D=0
M1 VSS A2 7 VSS N L=1.8e-07 W=1e-06 $X=1460 $Y=345 $D=0
M2 Z 6 VSS VSS N L=1.8e-07 W=1e-06 $X=2180 $Y=345 $D=0
M3 VSS 6 Z VSS N L=1.8e-07 W=1e-06 $X=2900 $Y=345 $D=0
M4 6 A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=740 $Y=2205 $D=16
M5 VDD A2 6 VDD P L=1.8e-07 W=1.37e-06 $X=1460 $Y=2205 $D=16
M6 Z 6 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2180 $Y=2205 $D=16
M7 VDD 6 Z VDD P L=1.8e-07 W=1.37e-06 $X=2900 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT IND2D2BWP7T A1 B1 ZN VSS VDD
** N=8 EP=5 IP=0 FDC=10
M0 VSS A1 6 VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 7 6 VSS VSS N L=1.8e-07 W=1e-06 $X=1420 $Y=345 $D=0
M2 ZN B1 7 VSS N L=1.8e-07 W=1e-06 $X=2060 $Y=345 $D=0
M3 8 B1 ZN VSS N L=1.8e-07 W=1e-06 $X=2780 $Y=345 $D=0
M4 VSS 6 8 VSS N L=1.8e-07 W=1e-06 $X=3380 $Y=345 $D=0
M5 VDD A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M6 ZN 6 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M7 VDD B1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M8 ZN B1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M9 VDD 6 ZN VDD P L=1.8e-07 W=1.37e-06 $X=3500 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300 301
+ 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321
+ 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341
+ 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361
+ 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381
+ 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401
+ 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421
+ 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441
+ 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461
+ 462 463 464 465 466 467 468 469 470 471 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696
** N=1302 EP=694 IP=6353 FDC=10288
M0 1 950 877 1 N L=1.8e-07 W=5e-07 $X=81100 $Y=263385 $D=0
M1 950 4 1294 1 N L=1.8e-07 W=5e-07 $X=82370 $Y=263760 $D=0
M2 1294 946 950 1 N L=1.8e-07 W=5e-07 $X=83090 $Y=263760 $D=0
M3 1295 909 1294 1 N L=1.8e-07 W=5e-07 $X=83690 $Y=263385 $D=0
M4 1 947 1295 1 N L=1.8e-07 W=5e-07 $X=84140 $Y=263385 $D=0
M5 1 241 1082 1 N L=1.8e-07 W=5e-07 $X=185820 $Y=238425 $D=0
M6 1296 1086 1 1 N L=1.8e-07 W=5e-07 $X=186580 $Y=238245 $D=0
M7 1096 241 1296 1 N L=1.8e-07 W=5e-07 $X=187160 $Y=238245 $D=0
M8 1086 1082 1096 1 N L=1.8e-07 W=5e-07 $X=187880 $Y=238245 $D=0
M9 1 1087 1086 1 N L=1.8e-07 W=1e-06 $X=188660 $Y=238175 $D=0
M10 254 1095 1 1 N L=1.8e-07 W=1e-06 $X=189420 $Y=238175 $D=0
M11 1 1095 254 1 N L=1.8e-07 W=1e-06 $X=190140 $Y=238175 $D=0
M12 1095 1098 1096 1 N L=1.8e-07 W=5e-07 $X=191570 $Y=238580 $D=0
M13 1297 1097 1095 1 N L=1.8e-07 W=5e-07 $X=192330 $Y=238175 $D=0
M14 1 1096 1297 1 N L=1.8e-07 W=5e-07 $X=192810 $Y=238175 $D=0
M15 1097 1098 1 1 N L=1.8e-07 W=5e-07 $X=193530 $Y=238175 $D=0
M16 1099 266 1 1 N L=1.8e-07 W=1e-06 $X=194950 $Y=238175 $D=0
M17 1098 1102 1099 1 N L=1.8e-07 W=5e-07 $X=195730 $Y=238245 $D=0
M18 1298 1100 1098 1 N L=1.8e-07 W=5e-07 $X=196450 $Y=238245 $D=0
M19 1 1099 1298 1 N L=1.8e-07 W=5e-07 $X=197080 $Y=238245 $D=0
M20 1102 1100 1 1 N L=1.8e-07 W=5e-07 $X=197840 $Y=238420 $D=0
M21 2 950 877 2 P L=1.8e-07 W=6.85e-07 $X=81315 $Y=265930 $D=16
M22 1299 4 2 2 P L=1.8e-07 W=6.85e-07 $X=82115 $Y=265930 $D=16
M23 950 946 1299 2 P L=1.8e-07 W=6.85e-07 $X=82695 $Y=265930 $D=16
M24 2 909 950 2 P L=1.8e-07 W=6.85e-07 $X=83415 $Y=265930 $D=16
M25 950 947 2 2 P L=1.8e-07 W=6.85e-07 $X=84140 $Y=265930 $D=16
M26 2 241 1082 2 P L=1.8e-07 W=6.85e-07 $X=185820 $Y=236115 $D=16
M27 1300 1086 2 2 P L=1.8e-07 W=6.85e-07 $X=186580 $Y=236450 $D=16
M28 1096 1082 1300 2 P L=1.8e-07 W=6.85e-07 $X=187160 $Y=236450 $D=16
M29 1086 241 1096 2 P L=1.8e-07 W=6.85e-07 $X=187880 $Y=236450 $D=16
M30 2 1087 1086 2 P L=1.8e-07 W=1.37e-06 $X=188660 $Y=235945 $D=16
M31 254 1095 2 2 P L=1.8e-07 W=1.37e-06 $X=189420 $Y=235945 $D=16
M32 2 1095 254 2 P L=1.8e-07 W=1.37e-06 $X=190140 $Y=235945 $D=16
M33 1095 1097 1096 2 P L=1.8e-07 W=6.85e-07 $X=191580 $Y=236430 $D=16
M34 1301 1098 1095 2 P L=1.8e-07 W=6.85e-07 $X=192320 $Y=236430 $D=16
M35 2 1096 1301 2 P L=1.8e-07 W=6.85e-07 $X=192810 $Y=236430 $D=16
M36 1097 1098 2 2 P L=1.8e-07 W=6.85e-07 $X=193530 $Y=236430 $D=16
M37 1099 266 2 2 P L=1.8e-07 W=1.37e-06 $X=194990 $Y=235945 $D=16
M38 1098 1100 1099 2 P L=1.8e-07 W=6.85e-07 $X=195710 $Y=236405 $D=16
M39 1302 1102 1098 2 P L=1.8e-07 W=6.85e-07 $X=196450 $Y=236405 $D=16
M40 2 1099 1302 2 P L=1.8e-07 W=6.85e-07 $X=197080 $Y=236405 $D=16
M41 1102 1100 2 2 P L=1.8e-07 W=6.85e-07 $X=197840 $Y=236160 $D=16
X111 1 674 ANTENNABWP7T $T=473040 231680 0 0 $X=472750 $Y=231445
X112 1 691 ANTENNABWP7T $T=474160 239520 0 180 $X=472750 $Y=235310
X113 1 690 ANTENNABWP7T $T=473040 239520 0 0 $X=472750 $Y=239285
X114 1 596 ANTENNABWP7T $T=474160 247360 0 180 $X=472750 $Y=243150
X115 1 561 ANTENNABWP7T $T=473040 247360 0 0 $X=472750 $Y=247125
X116 1 548 ANTENNABWP7T $T=474160 255200 0 180 $X=472750 $Y=250990
X117 1 411 ANTENNABWP7T $T=473040 255200 0 0 $X=472750 $Y=254965
X118 1 671 ANTENNABWP7T $T=473040 263040 0 0 $X=472750 $Y=262805
X119 1 678 ANTENNABWP7T $T=474160 270880 0 180 $X=472750 $Y=266670
X120 1 689 ANTENNABWP7T $T=473040 270880 0 0 $X=472750 $Y=270645
X121 1 692 ANTENNABWP7T $T=474160 278720 0 180 $X=472750 $Y=274510
X122 1 695 ANTENNABWP7T $T=473040 278720 0 0 $X=472750 $Y=278485
X123 1 693 ANTENNABWP7T $T=474160 286560 0 180 $X=472750 $Y=282350
X124 1 659 ANTENNABWP7T $T=473040 286560 0 0 $X=472750 $Y=286325
X125 1 582 675 ICV_1 $T=470800 231680 0 0 $X=470510 $Y=231445
X126 1 679 696 ICV_1 $T=470800 239520 0 0 $X=470510 $Y=239285
X127 1 672 683 ICV_1 $T=470800 247360 0 0 $X=470510 $Y=247125
X128 1 645 408 ICV_1 $T=470800 255200 0 0 $X=470510 $Y=254965
X129 1 680 684 ICV_1 $T=470800 263040 0 0 $X=470510 $Y=262805
X130 1 581 677 ICV_1 $T=470800 270880 0 0 $X=470510 $Y=270645
X131 1 461 685 ICV_1 $T=470800 278720 0 0 $X=470510 $Y=278485
X132 1 638 666 ICV_1 $T=470800 286560 0 0 $X=470510 $Y=286325
X133 1 487 617 ICV_2 $T=470800 263040 0 180 $X=469390 $Y=258830
X134 1 644 530 ICV_2 $T=471920 239520 0 180 $X=470510 $Y=235310
X135 1 657 673 ICV_2 $T=471920 247360 0 180 $X=470510 $Y=243150
X136 1 594 604 ICV_2 $T=471920 255200 0 180 $X=470510 $Y=250990
X137 1 609 668 ICV_2 $T=471920 270880 0 180 $X=470510 $Y=266670
X138 1 686 403 ICV_2 $T=471920 278720 0 180 $X=470510 $Y=274510
X139 1 687 682 ICV_2 $T=471920 286560 0 180 $X=470510 $Y=282350
X140 1 484 439 ICV_2 $T=473040 263040 0 180 $X=471630 $Y=258830
X141 1 694 688 ICV_2 $T=473040 294400 0 180 $X=471630 $Y=290190
X235 170 1 2 1017 CKBD1BWP7T $T=135920 239520 1 0 $X=135630 $Y=235310
X236 183 1 2 1024 CKBD1BWP7T $T=146000 278720 0 0 $X=145710 $Y=278485
X237 189 1 2 1034 CKBD1BWP7T $T=149360 294400 1 0 $X=149070 $Y=290190
X238 285 1 2 1104 CKBD1BWP7T $T=210960 278720 1 0 $X=210670 $Y=274510
X239 1114 1 2 295 CKBD1BWP7T $T=221040 278720 1 0 $X=220750 $Y=274510
X240 398 1 2 1176 CKBD1BWP7T $T=279840 294400 0 180 $X=277310 $Y=290190
X241 403 1 2 1171 CKBD1BWP7T $T=282080 255200 1 180 $X=279550 $Y=254965
X242 404 1 2 1180 CKBD1BWP7T $T=282080 294400 0 180 $X=279550 $Y=290190
X243 408 1 2 1169 CKBD1BWP7T $T=292160 263040 1 180 $X=289630 $Y=262805
X244 411 1 2 1177 CKBD1BWP7T $T=293280 247360 0 180 $X=290750 $Y=243150
X245 439 1 2 1192 CKBD1BWP7T $T=308400 255200 0 180 $X=305870 $Y=250990
X246 1198 1 2 1127 CKBD1BWP7T $T=308400 270880 1 180 $X=305870 $Y=270645
X247 469 1 2 471 CKBD1BWP7T $T=322960 270880 0 0 $X=322670 $Y=270645
X248 487 1 2 456 CKBD1BWP7T $T=342000 263040 1 180 $X=339470 $Y=262805
X249 591 1 2 640 CKBD1BWP7T $T=448960 270880 0 0 $X=448670 $Y=270645
X250 644 1 2 641 CKBD1BWP7T $T=460720 247360 1 180 $X=458190 $Y=247125
X251 650 1 2 1186 CKBD1BWP7T $T=462400 286560 0 180 $X=459870 $Y=282350
X252 881 1 2 857 INVD0BWP7T $T=45200 247360 0 180 $X=43230 $Y=243150
X253 935 1 2 939 INVD0BWP7T $T=71520 263040 1 0 $X=71230 $Y=258830
X254 927 1 2 936 INVD0BWP7T $T=71520 286560 0 0 $X=71230 $Y=286325
X255 107 1 2 114 INVD0BWP7T $T=93360 231680 0 0 $X=93070 $Y=231445
X256 954 1 2 103 INVD0BWP7T $T=96160 278720 0 0 $X=95870 $Y=278485
X257 984 1 2 976 INVD0BWP7T $T=109040 263040 0 180 $X=107070 $Y=258830
X258 890 1 2 971 INVD0BWP7T $T=107920 286560 1 0 $X=107630 $Y=282350
X259 983 1 2 982 INVD0BWP7T $T=110160 247360 1 180 $X=108190 $Y=247125
X260 54 1 2 994 INVD0BWP7T $T=121920 239520 0 0 $X=121630 $Y=239285
X261 62 1 2 1012 INVD0BWP7T $T=143760 270880 1 180 $X=141790 $Y=270645
X262 1005 1 2 175 INVD0BWP7T $T=143760 270880 0 0 $X=143470 $Y=270645
X263 1034 1 2 1039 INVD0BWP7T $T=151600 286560 1 0 $X=151310 $Y=282350
X264 176 1 2 1031 INVD0BWP7T $T=152160 270880 0 0 $X=151870 $Y=270645
X265 195 1 2 1026 INVD0BWP7T $T=153280 255200 0 0 $X=152990 $Y=254965
X266 210 1 2 1048 INVD0BWP7T $T=163920 239520 1 0 $X=163630 $Y=235310
X267 1049 1 2 1043 INVD0BWP7T $T=165600 239520 1 180 $X=163630 $Y=239285
X268 1032 1 2 1062 INVD0BWP7T $T=170640 278720 0 0 $X=170350 $Y=278485
X269 1059 1 2 1060 INVD0BWP7T $T=171200 270880 0 0 $X=170910 $Y=270645
X270 1037 1 2 1078 INVD0BWP7T $T=182960 255200 1 0 $X=182670 $Y=250990
X271 1061 1 2 1081 INVD0BWP7T $T=186320 270880 0 0 $X=186030 $Y=270645
X272 1137 1 2 1141 INVD0BWP7T $T=248480 239520 0 0 $X=248190 $Y=239285
X273 1150 1 2 1149 INVD0BWP7T $T=255760 239520 1 180 $X=253790 $Y=239285
X274 354 1 2 1158 INVD0BWP7T $T=261920 239520 1 0 $X=261630 $Y=235310
X275 382 1 2 1175 INVD0BWP7T $T=273120 278720 0 0 $X=272830 $Y=278485
X276 403 1 2 1168 INVD0BWP7T $T=291600 263040 0 180 $X=289630 $Y=258830
X277 408 1 2 1172 INVD0BWP7T $T=294960 255200 1 180 $X=292990 $Y=254965
X278 411 1 2 1181 INVD0BWP7T $T=301120 247360 0 180 $X=299150 $Y=243150
X279 439 1 2 1201 INVD0BWP7T $T=308960 255200 1 0 $X=308670 $Y=250990
X280 1209 1 2 1210 INVD0BWP7T $T=335280 247360 0 0 $X=334990 $Y=247125
X281 488 1 2 1216 INVD0BWP7T $T=340880 239520 1 0 $X=340590 $Y=235310
X282 484 1 2 1214 INVD0BWP7T $T=351520 263040 0 0 $X=351230 $Y=262805
X283 1227 1 2 1218 INVD0BWP7T $T=358240 286560 0 180 $X=356270 $Y=282350
X284 1228 1 2 1225 INVD0BWP7T $T=361040 263040 0 0 $X=360750 $Y=262805
X285 528 1 2 1236 INVD0BWP7T $T=378400 278720 1 180 $X=376430 $Y=278485
X286 524 1 2 1234 INVD0BWP7T $T=376720 286560 1 0 $X=376430 $Y=282350
X287 236 1 2 1231 INVD0BWP7T $T=377280 263040 0 0 $X=376990 $Y=262805
X288 534 1 2 1239 INVD0BWP7T $T=382320 263040 0 180 $X=380350 $Y=258830
X289 1246 1 2 1243 INVD0BWP7T $T=392400 286560 1 180 $X=390430 $Y=286325
X290 1247 1 2 558 INVD0BWP7T $T=398000 294400 0 180 $X=396030 $Y=290190
X291 1252 1 2 1256 INVD0BWP7T $T=406960 247360 1 0 $X=406670 $Y=243150
X292 576 1 2 1261 INVD0BWP7T $T=417600 286560 1 0 $X=417310 $Y=282350
X293 1265 1 2 593 INVD0BWP7T $T=422640 294400 1 0 $X=422350 $Y=290190
X294 547 1 2 605 INVD0BWP7T $T=432160 231680 0 0 $X=431870 $Y=231445
X295 272 1 2 1271 INVD0BWP7T $T=438880 255200 1 0 $X=438590 $Y=250990
X296 635 1 2 1269 INVD0BWP7T $T=446720 239520 0 180 $X=444750 $Y=235310
X297 582 1 2 1274 INVD0BWP7T $T=448400 239520 1 0 $X=448110 $Y=235310
X298 624 1 2 632 INVD0BWP7T $T=450640 231680 1 180 $X=448670 $Y=231445
X299 1162 1 2 1277 INVD0BWP7T $T=457920 263040 1 0 $X=457630 $Y=258830
X300 643 1 2 1275 INVD0BWP7T $T=459600 247360 1 0 $X=459310 $Y=243150
X301 649 1 2 1278 INVD0BWP7T $T=460720 247360 0 0 $X=460430 $Y=247125
X302 508 1 2 1276 INVD0BWP7T $T=462960 247360 0 180 $X=460990 $Y=243150
X303 317 1 2 1280 INVD0BWP7T $T=461280 278720 0 0 $X=460990 $Y=278485
X304 654 1 2 1279 INVD0BWP7T $T=464080 263040 0 180 $X=462110 $Y=258830
X305 656 1 2 1281 INVD0BWP7T $T=462960 270880 0 0 $X=462670 $Y=270645
X306 995 203 1 2 BUFFD1P5BWP7T $T=153280 239520 0 0 $X=152990 $Y=239285
X307 1058 245 1 2 BUFFD1P5BWP7T $T=179040 231680 0 0 $X=178750 $Y=231445
X308 276 284 1 2 BUFFD1P5BWP7T $T=207040 286560 1 0 $X=206750 $Y=282350
X309 1138 334 1 2 BUFFD1P5BWP7T $T=247920 270880 1 0 $X=247630 $Y=266670
X310 1093 416 1 2 BUFFD1P5BWP7T $T=291600 263040 1 0 $X=291310 $Y=258830
X311 461 392 1 2 BUFFD1P5BWP7T $T=320160 286560 0 180 $X=317070 $Y=282350
X312 1092 489 1 2 BUFFD1P5BWP7T $T=340320 270880 0 0 $X=340030 $Y=270645
X313 530 526 1 2 BUFFD1P5BWP7T $T=379520 239520 1 180 $X=376430 $Y=239285
X314 548 546 1 2 BUFFD1P5BWP7T $T=391840 263040 0 180 $X=388750 $Y=258830
X315 561 560 1 2 BUFFD1P5BWP7T $T=400240 247360 0 180 $X=397150 $Y=243150
X316 581 583 1 2 BUFFD1P5BWP7T $T=417040 270880 0 0 $X=416750 $Y=270645
X317 594 458 1 2 BUFFD1P5BWP7T $T=425440 247360 1 180 $X=422350 $Y=247125
X318 596 572 1 2 BUFFD1P5BWP7T $T=426000 247360 0 180 $X=422910 $Y=243150
X319 1266 601 1 2 BUFFD1P5BWP7T $T=426560 255200 0 0 $X=426270 $Y=254965
X320 602 598 1 2 BUFFD1P5BWP7T $T=429920 294400 0 180 $X=426830 $Y=290190
X321 604 462 1 2 BUFFD1P5BWP7T $T=431600 247360 0 180 $X=428510 $Y=243150
X322 609 589 1 2 BUFFD1P5BWP7T $T=435520 263040 1 180 $X=432430 $Y=262805
X323 617 614 1 2 BUFFD1P5BWP7T $T=438880 239520 1 180 $X=435790 $Y=239285
X324 645 1128 1 2 BUFFD1P5BWP7T $T=460720 255200 1 180 $X=457630 $Y=254965
X325 648 642 1 2 BUFFD1P5BWP7T $T=461840 270880 0 180 $X=458750 $Y=266670
X326 651 646 1 2 BUFFD1P5BWP7T $T=462400 286560 1 180 $X=459310 $Y=286325
X327 652 532 1 2 BUFFD1P5BWP7T $T=462960 294400 0 180 $X=459870 $Y=290190
X328 657 528 1 2 BUFFD1P5BWP7T $T=464640 270880 0 180 $X=461550 $Y=266670
X329 659 655 1 2 BUFFD1P5BWP7T $T=465760 294400 0 180 $X=462670 $Y=290190
X330 666 348 1 2 BUFFD1P5BWP7T $T=469120 286560 0 180 $X=466030 $Y=282350
X331 668 622 1 2 BUFFD1P5BWP7T $T=469680 263040 0 180 $X=466590 $Y=258830
X332 672 670 1 2 BUFFD1P5BWP7T $T=470800 239520 0 180 $X=467710 $Y=235310
X333 673 667 1 2 BUFFD1P5BWP7T $T=470800 239520 1 180 $X=467710 $Y=239285
X334 674 1162 1 2 BUFFD1P5BWP7T $T=470800 247360 1 180 $X=467710 $Y=247125
X335 675 664 1 2 BUFFD1P5BWP7T $T=470800 278720 0 180 $X=467710 $Y=274510
X336 676 665 1 2 BUFFD1P5BWP7T $T=470800 278720 1 180 $X=467710 $Y=278485
X337 677 478 1 2 BUFFD1P5BWP7T $T=470800 286560 1 180 $X=467710 $Y=286325
X338 669 1 2 681 INVD3BWP7T $T=468560 294400 1 0 $X=468270 $Y=290190
X339 1168 388 2 1 388 1173 1168 MAOI22D0BWP7T $T=279280 255200 0 180 $X=275070 $Y=250990
X340 392 1176 2 1 392 1179 1180 MAOI22D0BWP7T $T=277040 286560 0 0 $X=276750 $Y=286325
X341 1172 415 2 1 415 1178 1172 MAOI22D0BWP7T $T=296080 255200 0 180 $X=291870 $Y=250990
X342 440 428 2 1 440 1200 428 MAOI22D0BWP7T $T=312320 278720 1 180 $X=308110 $Y=278485
X343 598 1257 2 1 598 597 1257 MAOI22D0BWP7T $T=430480 231680 1 180 $X=426270 $Y=231445
X412 258 205 205 258 1087 1 2 MAOI22D2BWP7T $T=193040 263040 0 0 $X=192750 $Y=262805
X413 622 619 622 619 616 1 2 MAOI22D2BWP7T $T=442800 239520 0 180 $X=436350 $Y=235310
X414 661 660 661 660 1184 1 2 MAOI22D2BWP7T $T=469120 263040 1 180 $X=462670 $Y=262805
X415 213 210 204 213 1 210 2 IAO22D2BWP7T $T=170080 255200 0 180 $X=163630 $Y=250990
X416 572 586 577 572 1 586 2 IAO22D2BWP7T $T=426560 270880 0 180 $X=420110 $Y=266670
X417 866 1 2 30 BUFFD1BWP7T $T=39040 294400 1 0 $X=38750 $Y=290190
X418 60 1 2 905 BUFFD1BWP7T $T=59760 239520 0 180 $X=57230 $Y=235310
X419 911 1 2 79 BUFFD1BWP7T $T=65920 255200 0 0 $X=65630 $Y=254965
X420 942 1 2 945 BUFFD1BWP7T $T=79920 270880 0 0 $X=79630 $Y=270645
X421 956 1 2 138 BUFFD1BWP7T $T=107360 231680 0 0 $X=107070 $Y=231445
X422 1003 1 2 1008 BUFFD1BWP7T $T=126960 231680 0 0 $X=126670 $Y=231445
X423 173 1 2 1018 BUFFD1BWP7T $T=138160 239520 1 0 $X=137870 $Y=235310
X424 930 1 2 1022 BUFFD1BWP7T $T=142640 286560 0 0 $X=142350 $Y=286325
X425 1025 1 2 1032 BUFFD1BWP7T $T=148240 278720 0 0 $X=147950 $Y=278485
X426 1009 1 2 207 BUFFD1BWP7T $T=154960 255200 0 0 $X=154670 $Y=254965
X427 294 1 2 1115 BUFFD1BWP7T $T=220480 278720 0 0 $X=220190 $Y=278485
X428 1161 1 2 1144 BUFFD1BWP7T $T=262480 255200 1 180 $X=259950 $Y=254965
X429 377 1 2 374 BUFFD1BWP7T $T=271440 286560 1 180 $X=268910 $Y=286325
X430 1094 1 2 410 BUFFD1BWP7T $T=289920 270880 1 0 $X=289630 $Y=266670
X431 1203 1 2 455 BUFFD1BWP7T $T=320160 270880 0 180 $X=317630 $Y=266670
X432 1205 1 2 467 BUFFD1BWP7T $T=319600 278720 0 0 $X=319310 $Y=278485
X433 1204 1 2 466 BUFFD1BWP7T $T=320160 270880 1 0 $X=319870 $Y=266670
X434 1225 1 2 1224 BUFFD1BWP7T $T=357680 263040 0 0 $X=357390 $Y=262805
X435 1226 1 2 1229 BUFFD1BWP7T $T=361040 255200 1 0 $X=360750 $Y=250990
X436 562 1 2 565 BUFFD1BWP7T $T=406960 255200 0 0 $X=406670 $Y=254965
X437 1270 1 2 637 BUFFD1BWP7T $T=445040 255200 1 0 $X=444750 $Y=250990
X438 1272 1 2 653 BUFFD1BWP7T $T=457920 231680 0 0 $X=457630 $Y=231445
X439 1 2 DCAP4BWP7T $T=21120 247360 1 0 $X=20830 $Y=243150
X440 1 2 DCAP4BWP7T $T=55280 255200 0 0 $X=54990 $Y=254965
X441 1 2 DCAP4BWP7T $T=64240 278720 1 0 $X=63950 $Y=274510
X442 1 2 DCAP4BWP7T $T=83280 278720 1 0 $X=82990 $Y=274510
X443 1 2 DCAP4BWP7T $T=101760 286560 0 0 $X=101470 $Y=286325
X444 1 2 DCAP4BWP7T $T=124160 270880 0 0 $X=123870 $Y=270645
X445 1 2 DCAP4BWP7T $T=145440 270880 0 0 $X=145150 $Y=270645
X446 1 2 DCAP4BWP7T $T=157760 263040 0 0 $X=157470 $Y=262805
X447 1 2 DCAP4BWP7T $T=182960 239520 0 0 $X=182670 $Y=239285
X448 1 2 DCAP4BWP7T $T=231120 247360 1 0 $X=230830 $Y=243150
X449 1 2 DCAP4BWP7T $T=283760 255200 1 0 $X=283470 $Y=250990
X450 1 2 DCAP4BWP7T $T=283760 263040 0 0 $X=283470 $Y=262805
X451 1 2 DCAP4BWP7T $T=301120 247360 1 0 $X=300830 $Y=243150
X452 1 2 DCAP4BWP7T $T=303920 255200 1 0 $X=303630 $Y=250990
X453 1 2 DCAP4BWP7T $T=338080 270880 0 0 $X=337790 $Y=270645
X454 1 2 DCAP4BWP7T $T=349280 247360 0 0 $X=348990 $Y=247125
X455 1 2 DCAP4BWP7T $T=367760 231680 0 0 $X=367470 $Y=231445
X456 1 2 DCAP4BWP7T $T=367760 255200 1 0 $X=367470 $Y=250990
X457 1 2 DCAP4BWP7T $T=435520 270880 1 0 $X=435230 $Y=266670
X458 1 2 DCAP4BWP7T $T=451760 278720 1 0 $X=451470 $Y=274510
X459 1 2 DCAP4BWP7T $T=465760 239520 1 0 $X=465470 $Y=235310
X460 1 2 ICV_3 $T=31200 255200 0 0 $X=30910 $Y=254965
X461 1 2 ICV_3 $T=31200 263040 1 0 $X=30910 $Y=258830
X462 1 2 ICV_3 $T=31200 270880 1 0 $X=30910 $Y=266670
X463 1 2 ICV_3 $T=31200 278720 0 0 $X=30910 $Y=278485
X464 1 2 ICV_3 $T=31200 294400 1 0 $X=30910 $Y=290190
X465 1 2 ICV_3 $T=35120 286560 0 0 $X=34830 $Y=286325
X466 1 2 ICV_3 $T=54160 239520 0 0 $X=53870 $Y=239285
X467 1 2 ICV_3 $T=86640 294400 1 0 $X=86350 $Y=290190
X468 1 2 ICV_3 $T=109600 286560 1 0 $X=109310 $Y=282350
X469 1 2 ICV_3 $T=115200 278720 0 0 $X=114910 $Y=278485
X470 1 2 ICV_3 $T=115200 294400 1 0 $X=114910 $Y=290190
X471 1 2 ICV_3 $T=119120 255200 0 0 $X=118830 $Y=254965
X472 1 2 ICV_3 $T=146000 231680 0 0 $X=145710 $Y=231445
X473 1 2 ICV_3 $T=157200 231680 0 0 $X=156910 $Y=231445
X474 1 2 ICV_3 $T=157200 239520 1 0 $X=156910 $Y=235310
X475 1 2 ICV_3 $T=157200 247360 1 0 $X=156910 $Y=243150
X476 1 2 ICV_3 $T=157200 255200 0 0 $X=156910 $Y=254965
X477 1 2 ICV_3 $T=157200 263040 1 0 $X=156910 $Y=258830
X478 1 2 ICV_3 $T=157200 270880 1 0 $X=156910 $Y=266670
X479 1 2 ICV_3 $T=157200 278720 1 0 $X=156910 $Y=274510
X480 1 2 ICV_3 $T=157200 278720 0 0 $X=156910 $Y=278485
X481 1 2 ICV_3 $T=157200 294400 1 0 $X=156910 $Y=290190
X482 1 2 ICV_3 $T=183520 263040 1 0 $X=183230 $Y=258830
X483 1 2 ICV_3 $T=199200 247360 0 0 $X=198910 $Y=247125
X484 1 2 ICV_3 $T=199200 255200 0 0 $X=198910 $Y=254965
X485 1 2 ICV_3 $T=199200 263040 0 0 $X=198910 $Y=262805
X486 1 2 ICV_3 $T=199200 270880 1 0 $X=198910 $Y=266670
X487 1 2 ICV_3 $T=199200 278720 1 0 $X=198910 $Y=274510
X488 1 2 ICV_3 $T=199200 278720 0 0 $X=198910 $Y=278485
X489 1 2 ICV_3 $T=203120 270880 0 0 $X=202830 $Y=270645
X490 1 2 ICV_3 $T=231120 294400 1 0 $X=230830 $Y=290190
X491 1 2 ICV_3 $T=241200 239520 1 0 $X=240910 $Y=235310
X492 1 2 ICV_3 $T=245120 270880 1 0 $X=244830 $Y=266670
X493 1 2 ICV_3 $T=264720 255200 1 0 $X=264430 $Y=250990
X494 1 2 ICV_3 $T=291600 247360 0 0 $X=291310 $Y=247125
X495 1 2 ICV_3 $T=301680 286560 1 0 $X=301390 $Y=282350
X496 1 2 ICV_3 $T=306160 270880 1 0 $X=305870 $Y=266670
X497 1 2 ICV_3 $T=315120 255200 1 0 $X=314830 $Y=250990
X498 1 2 ICV_3 $T=316800 278720 0 0 $X=316510 $Y=278485
X499 1 2 ICV_3 $T=333600 263040 1 0 $X=333310 $Y=258830
X500 1 2 ICV_3 $T=409200 231680 0 0 $X=408910 $Y=231445
X501 1 2 ICV_3 $T=409200 255200 0 0 $X=408910 $Y=254965
X502 1 2 ICV_3 $T=424320 294400 1 0 $X=424030 $Y=290190
X503 1 2 ICV_3 $T=426000 247360 1 0 $X=425710 $Y=243150
X504 1 2 ICV_3 $T=446160 231680 0 0 $X=445870 $Y=231445
X505 1 2 ICV_3 $T=446160 270880 0 0 $X=445870 $Y=270645
X506 1 2 ICV_3 $T=464080 263040 1 0 $X=463790 $Y=258830
X507 1 2 ICV_3 $T=464640 270880 1 0 $X=464350 $Y=266670
X508 1 2 ICV_3 $T=465760 294400 1 0 $X=465470 $Y=290190
X509 1 2 DCAP8BWP7T $T=27840 263040 0 0 $X=27550 $Y=262805
X510 1 2 DCAP8BWP7T $T=27840 278720 1 0 $X=27550 $Y=274510
X511 1 2 DCAP8BWP7T $T=28960 239520 0 0 $X=28670 $Y=239285
X512 1 2 DCAP8BWP7T $T=52480 270880 0 0 $X=52190 $Y=270645
X513 1 2 DCAP8BWP7T $T=53040 247360 1 0 $X=52750 $Y=243150
X514 1 2 DCAP8BWP7T $T=56960 247360 0 0 $X=56670 $Y=247125
X515 1 2 DCAP8BWP7T $T=57520 231680 0 0 $X=57230 $Y=231445
X516 1 2 DCAP8BWP7T $T=66480 263040 1 0 $X=66190 $Y=258830
X517 1 2 DCAP8BWP7T $T=70960 239520 1 0 $X=70670 $Y=235310
X518 1 2 DCAP8BWP7T $T=93920 263040 1 0 $X=93630 $Y=258830
X519 1 2 DCAP8BWP7T $T=119120 231680 0 0 $X=118830 $Y=231445
X520 1 2 DCAP8BWP7T $T=128080 247360 1 0 $X=127790 $Y=243150
X521 1 2 DCAP8BWP7T $T=129200 247360 0 0 $X=128910 $Y=247125
X522 1 2 DCAP8BWP7T $T=130320 270880 0 0 $X=130030 $Y=270645
X523 1 2 DCAP8BWP7T $T=133680 270880 1 0 $X=133390 $Y=266670
X524 1 2 DCAP8BWP7T $T=144320 294400 1 0 $X=144030 $Y=290190
X525 1 2 DCAP8BWP7T $T=161120 286560 1 0 $X=160830 $Y=282350
X526 1 2 DCAP8BWP7T $T=197520 231680 0 0 $X=197230 $Y=231445
X527 1 2 DCAP8BWP7T $T=197520 247360 1 0 $X=197230 $Y=243150
X528 1 2 DCAP8BWP7T $T=197520 286560 0 0 $X=197230 $Y=286325
X529 1 2 DCAP8BWP7T $T=214320 286560 0 0 $X=214030 $Y=286325
X530 1 2 DCAP8BWP7T $T=217680 255200 0 0 $X=217390 $Y=254965
X531 1 2 DCAP8BWP7T $T=218240 263040 1 0 $X=217950 $Y=258830
X532 1 2 DCAP8BWP7T $T=220480 247360 1 0 $X=220190 $Y=243150
X533 1 2 DCAP8BWP7T $T=237840 247360 0 0 $X=237550 $Y=247125
X534 1 2 DCAP8BWP7T $T=239520 239520 0 0 $X=239230 $Y=239285
X535 1 2 DCAP8BWP7T $T=239520 247360 1 0 $X=239230 $Y=243150
X536 1 2 DCAP8BWP7T $T=239520 270880 0 0 $X=239230 $Y=270645
X537 1 2 DCAP8BWP7T $T=245120 255200 0 0 $X=244830 $Y=254965
X538 1 2 DCAP8BWP7T $T=250720 270880 1 0 $X=250430 $Y=266670
X539 1 2 DCAP8BWP7T $T=255760 286560 1 0 $X=255470 $Y=282350
X540 1 2 DCAP8BWP7T $T=263600 239520 1 0 $X=263310 $Y=235310
X541 1 2 DCAP8BWP7T $T=266400 278720 1 0 $X=266110 $Y=274510
X542 1 2 DCAP8BWP7T $T=270320 286560 1 0 $X=270030 $Y=282350
X543 1 2 DCAP8BWP7T $T=279840 286560 1 0 $X=279550 $Y=282350
X544 1 2 DCAP8BWP7T $T=280960 286560 0 0 $X=280670 $Y=286325
X545 1 2 DCAP8BWP7T $T=294400 263040 1 0 $X=294110 $Y=258830
X546 1 2 DCAP8BWP7T $T=323520 239520 0 0 $X=323230 $Y=239285
X547 1 2 DCAP8BWP7T $T=329120 294400 1 0 $X=328830 $Y=290190
X548 1 2 DCAP8BWP7T $T=334720 270880 1 0 $X=334430 $Y=266670
X549 1 2 DCAP8BWP7T $T=342000 239520 0 0 $X=341710 $Y=239285
X550 1 2 DCAP8BWP7T $T=342000 286560 1 0 $X=341710 $Y=282350
X551 1 2 DCAP8BWP7T $T=348720 294400 1 0 $X=348430 $Y=290190
X552 1 2 DCAP8BWP7T $T=353200 263040 0 0 $X=352910 $Y=262805
X553 1 2 DCAP8BWP7T $T=358240 286560 1 0 $X=357950 $Y=282350
X554 1 2 DCAP8BWP7T $T=364960 278720 1 0 $X=364670 $Y=274510
X555 1 2 DCAP8BWP7T $T=364960 286560 1 0 $X=364670 $Y=282350
X556 1 2 DCAP8BWP7T $T=365520 239520 1 0 $X=365230 $Y=235310
X557 1 2 DCAP8BWP7T $T=371120 278720 1 0 $X=370830 $Y=274510
X558 1 2 DCAP8BWP7T $T=382880 255200 0 0 $X=382590 $Y=254965
X559 1 2 DCAP8BWP7T $T=391840 263040 1 0 $X=391550 $Y=258830
X560 1 2 DCAP8BWP7T $T=395760 239520 0 0 $X=395470 $Y=239285
X561 1 2 DCAP8BWP7T $T=400800 255200 0 0 $X=400510 $Y=254965
X562 1 2 DCAP8BWP7T $T=420400 231680 0 0 $X=420110 $Y=231445
X563 1 2 DCAP8BWP7T $T=434400 270880 0 0 $X=434110 $Y=270645
X564 1 2 DCAP8BWP7T $T=438880 239520 0 0 $X=438590 $Y=239285
X565 1 2 DCAP8BWP7T $T=439440 294400 1 0 $X=439150 $Y=290190
X566 1 2 DCAP8BWP7T $T=448960 255200 0 0 $X=448670 $Y=254965
X567 2 1 DCAPBWP7T $T=21120 255200 1 0 $X=20830 $Y=250990
X568 2 1 DCAPBWP7T $T=21120 255200 0 0 $X=20830 $Y=254965
X569 2 1 DCAPBWP7T $T=32320 263040 0 0 $X=32030 $Y=262805
X570 2 1 DCAPBWP7T $T=32320 278720 1 0 $X=32030 $Y=274510
X571 2 1 DCAPBWP7T $T=41840 247360 1 0 $X=41550 $Y=243150
X572 2 1 DCAPBWP7T $T=41840 255200 0 0 $X=41550 $Y=254965
X573 2 1 DCAPBWP7T $T=43520 263040 0 0 $X=43230 $Y=262805
X574 2 1 DCAPBWP7T $T=46320 294400 1 0 $X=46030 $Y=290190
X575 2 1 DCAPBWP7T $T=48560 278720 0 0 $X=48270 $Y=278485
X576 2 1 DCAPBWP7T $T=60880 255200 0 0 $X=60590 $Y=254965
X577 2 1 DCAPBWP7T $T=62000 231680 0 0 $X=61710 $Y=231445
X578 2 1 DCAPBWP7T $T=64240 239520 1 0 $X=63950 $Y=235310
X579 2 1 DCAPBWP7T $T=99520 239520 1 0 $X=99230 $Y=235310
X580 2 1 DCAPBWP7T $T=105120 239520 0 0 $X=104830 $Y=239285
X581 2 1 DCAPBWP7T $T=142640 247360 1 0 $X=142350 $Y=243150
X582 2 1 DCAPBWP7T $T=142640 270880 1 0 $X=142350 $Y=266670
X583 2 1 DCAPBWP7T $T=158320 270880 0 0 $X=158030 $Y=270645
X584 2 1 DCAPBWP7T $T=165600 286560 1 0 $X=165310 $Y=282350
X585 2 1 DCAPBWP7T $T=165600 294400 1 0 $X=165310 $Y=290190
X586 2 1 DCAPBWP7T $T=177920 247360 1 0 $X=177630 $Y=243150
X587 2 1 DCAPBWP7T $T=200320 263040 1 0 $X=200030 $Y=258830
X588 2 1 DCAPBWP7T $T=218240 239520 0 0 $X=217950 $Y=239285
X589 2 1 DCAPBWP7T $T=218800 286560 0 0 $X=218510 $Y=286325
X590 2 1 DCAPBWP7T $T=220480 270880 1 0 $X=220190 $Y=266670
X591 2 1 DCAPBWP7T $T=221600 247360 0 0 $X=221310 $Y=247125
X592 2 1 DCAPBWP7T $T=226640 239520 1 0 $X=226350 $Y=235310
X593 2 1 DCAPBWP7T $T=227200 239520 0 0 $X=226910 $Y=239285
X594 2 1 DCAPBWP7T $T=232240 255200 1 0 $X=231950 $Y=250990
X595 2 1 DCAPBWP7T $T=242320 247360 0 0 $X=242030 $Y=247125
X596 2 1 DCAPBWP7T $T=242320 286560 0 0 $X=242030 $Y=286325
X597 2 1 DCAPBWP7T $T=249600 255200 0 0 $X=249310 $Y=254965
X598 2 1 DCAPBWP7T $T=259120 247360 1 0 $X=258830 $Y=243150
X599 2 1 DCAPBWP7T $T=259680 278720 1 0 $X=259390 $Y=274510
X600 2 1 DCAPBWP7T $T=260240 286560 1 0 $X=259950 $Y=282350
X601 2 1 DCAPBWP7T $T=263600 263040 1 0 $X=263310 $Y=258830
X602 2 1 DCAPBWP7T $T=274240 247360 1 0 $X=273950 $Y=243150
X603 2 1 DCAPBWP7T $T=276480 239520 1 0 $X=276190 $Y=235310
X604 2 1 DCAPBWP7T $T=284320 286560 1 0 $X=284030 $Y=282350
X605 2 1 DCAPBWP7T $T=312880 247360 1 0 $X=312590 $Y=243150
X606 2 1 DCAPBWP7T $T=326320 278720 0 0 $X=326030 $Y=278485
X607 2 1 DCAPBWP7T $T=333600 286560 1 0 $X=333310 $Y=282350
X608 2 1 DCAPBWP7T $T=335840 286560 0 0 $X=335550 $Y=286325
X609 2 1 DCAPBWP7T $T=344800 278720 0 0 $X=344510 $Y=278485
X610 2 1 DCAPBWP7T $T=345920 255200 0 0 $X=345630 $Y=254965
X611 2 1 DCAPBWP7T $T=353200 294400 1 0 $X=352910 $Y=290190
X612 2 1 DCAPBWP7T $T=368320 270880 1 0 $X=368030 $Y=266670
X613 2 1 DCAPBWP7T $T=368320 278720 0 0 $X=368030 $Y=278485
X614 2 1 DCAPBWP7T $T=375600 263040 0 0 $X=375310 $Y=262805
X615 2 1 DCAPBWP7T $T=402480 270880 0 0 $X=402190 $Y=270645
X616 2 1 DCAPBWP7T $T=405280 255200 0 0 $X=404990 $Y=254965
X617 2 1 DCAPBWP7T $T=410320 247360 0 0 $X=410030 $Y=247125
X618 2 1 DCAPBWP7T $T=410320 270880 0 0 $X=410030 $Y=270645
X619 2 1 DCAPBWP7T $T=410320 278720 0 0 $X=410030 $Y=278485
X620 2 1 DCAPBWP7T $T=419840 278720 1 0 $X=419550 $Y=274510
X621 2 1 DCAPBWP7T $T=419840 286560 0 0 $X=419550 $Y=286325
X622 2 1 DCAPBWP7T $T=446720 239520 1 0 $X=446430 $Y=235310
X623 2 1 DCAPBWP7T $T=452320 239520 1 0 $X=452030 $Y=235310
X624 2 1 DCAPBWP7T $T=452320 247360 1 0 $X=452030 $Y=243150
X625 2 1 DCAPBWP7T $T=459600 278720 0 0 $X=459310 $Y=278485
X626 2 1 DCAPBWP7T $T=469120 231680 0 0 $X=468830 $Y=231445
X627 2 1 DCAPBWP7T $T=469120 270880 0 0 $X=468830 $Y=270645
X628 2 1 DCAPBWP7T $T=469120 286560 1 0 $X=468830 $Y=282350
X629 301 304 306 305 302 274 1 2 1118 AO222D0BWP7T $T=229440 278720 1 180 $X=222990 $Y=278485
X630 301 275 300 1117 272 274 1 2 1119 AO222D0BWP7T $T=223840 255200 1 0 $X=223550 $Y=250990
X631 301 304 296 293 261 274 1 2 311 AO222D0BWP7T $T=225520 263040 0 0 $X=225230 $Y=262805
X632 301 326 1130 308 314 274 1 2 1120 AO222D0BWP7T $T=239520 247360 0 180 $X=233070 $Y=243150
X633 304 301 1127 1129 317 274 1 2 1122 AO222D0BWP7T $T=240640 278720 1 180 $X=234190 $Y=278485
X634 301 304 1117 1132 319 274 1 2 1125 AO222D0BWP7T $T=241200 270880 0 180 $X=234750 $Y=266670
X635 301 304 295 1143 335 274 1 2 1126 AO222D0BWP7T $T=254640 278720 1 180 $X=248190 $Y=278485
X636 301 304 343 339 280 274 1 2 332 AO222D0BWP7T $T=255760 286560 1 180 $X=249310 $Y=286325
X637 301 304 337 343 345 274 1 2 352 AO222D0BWP7T $T=250720 294400 1 0 $X=250430 $Y=290190
X638 348 395 400 391 394 381 1 2 1124 AO222D0BWP7T $T=281520 278720 1 180 $X=275070 $Y=278485
X639 1162 274 401 391 302 381 1 2 1154 AO222D0BWP7T $T=282080 263040 0 180 $X=275630 $Y=258830
X640 338 395 419 391 410 381 1 2 1183 AO222D0BWP7T $T=298880 270880 1 180 $X=292430 $Y=270645
X641 409 274 426 391 240 381 1 2 1187 AO222D0BWP7T $T=301680 270880 0 180 $X=295230 $Y=266670
X642 460 395 453 450 416 448 1 2 442 AO222D0BWP7T $T=319600 270880 1 180 $X=313150 $Y=270645
X643 301 304 1127 1199 454 451 1 2 1206 AO222D0BWP7T $T=314560 247360 1 0 $X=314270 $Y=243150
X644 444 395 475 450 256 448 1 2 490 AO222D0BWP7T $T=331920 278720 0 0 $X=331630 $Y=278485
X645 301 304 1199 485 436 451 1 2 1215 AO222D0BWP7T $T=335840 239520 0 0 $X=335550 $Y=239285
X646 304 513 511 339 508 451 1 2 1219 AO222D0BWP7T $T=362720 239520 1 180 $X=356270 $Y=239285
X647 513 326 553 542 310 451 1 2 1240 AO222D0BWP7T $T=395760 239520 1 180 $X=389310 $Y=239285
X648 513 326 554 551 550 549 1 2 1242 AO222D0BWP7T $T=395760 270880 1 180 $X=389310 $Y=270645
X649 304 513 559 1233 557 451 1 2 1241 AO222D0BWP7T $T=398560 239520 0 180 $X=392110 $Y=235310
X650 513 326 542 1250 564 451 1 2 1248 AO222D0BWP7T $T=395760 263040 0 0 $X=395470 $Y=262805
X651 513 326 1251 554 565 549 1 2 1244 AO222D0BWP7T $T=397440 270880 1 0 $X=397150 $Y=266670
X652 630 549 625 450 224 448 1 2 1268 AO222D0BWP7T $T=444480 247360 1 180 $X=438030 $Y=247125
X653 628 549 626 450 633 448 1 2 1273 AO222D0BWP7T $T=441120 263040 0 0 $X=440830 $Y=262805
X654 623 1 624 627 632 2 1272 634 OAI221D1BWP7T $T=441120 231680 0 0 $X=440830 $Y=231445
X655 623 1 272 635 1271 2 1270 1269 OAI221D1BWP7T $T=448400 239520 1 180 $X=443070 $Y=239285
X656 1 2 ICV_4 $T=35120 263040 1 0 $X=34830 $Y=258830
X657 1 2 ICV_4 $T=35120 294400 1 0 $X=34830 $Y=290190
X658 1 2 ICV_4 $T=47440 247360 1 0 $X=47150 $Y=243150
X659 1 2 ICV_4 $T=114080 247360 0 0 $X=113790 $Y=247125
X660 1 2 ICV_4 $T=114080 263040 0 0 $X=113790 $Y=262805
X661 1 2 ICV_4 $T=114080 270880 0 0 $X=113790 $Y=270645
X662 1 2 ICV_4 $T=128080 270880 1 0 $X=127790 $Y=266670
X663 1 2 ICV_4 $T=138160 270880 0 0 $X=137870 $Y=270645
X664 1 2 ICV_4 $T=149360 278720 1 0 $X=149070 $Y=274510
X665 1 2 ICV_4 $T=156080 239520 0 0 $X=155790 $Y=239285
X666 1 2 ICV_4 $T=156080 286560 0 0 $X=155790 $Y=286325
X667 1 2 ICV_4 $T=168960 231680 0 0 $X=168670 $Y=231445
X668 1 2 ICV_4 $T=198080 255200 1 0 $X=197790 $Y=250990
X669 1 2 ICV_4 $T=203120 278720 0 0 $X=202830 $Y=278485
X670 1 2 ICV_4 $T=203120 286560 1 0 $X=202830 $Y=282350
X671 1 2 ICV_4 $T=210960 270880 0 0 $X=210670 $Y=270645
X672 1 2 ICV_4 $T=240080 286560 1 0 $X=239790 $Y=282350
X673 1 2 ICV_4 $T=245120 263040 1 0 $X=244830 $Y=258830
X674 1 2 ICV_4 $T=282080 255200 0 0 $X=281790 $Y=254965
X675 1 2 ICV_4 $T=282080 270880 1 0 $X=281790 $Y=266670
X676 1 2 ICV_4 $T=282080 294400 1 0 $X=281790 $Y=290190
X677 1 2 ICV_4 $T=287120 239520 0 0 $X=286830 $Y=239285
X678 1 2 ICV_4 $T=314000 270880 1 0 $X=313710 $Y=266670
X679 1 2 ICV_4 $T=324080 263040 0 0 $X=323790 $Y=262805
X680 1 2 ICV_4 $T=324080 286560 0 0 $X=323790 $Y=286325
X681 1 2 ICV_4 $T=329120 231680 0 0 $X=328830 $Y=231445
X682 1 2 ICV_4 $T=329120 270880 1 0 $X=328830 $Y=266670
X683 1 2 ICV_4 $T=352080 286560 0 0 $X=351790 $Y=286325
X684 1 2 ICV_4 $T=366080 247360 0 0 $X=365790 $Y=247125
X685 1 2 ICV_4 $T=366080 286560 0 0 $X=365790 $Y=286325
X686 1 2 ICV_4 $T=383440 270880 1 0 $X=383150 $Y=266670
X687 1 2 ICV_4 $T=413120 231680 0 0 $X=412830 $Y=231445
X688 1 2 ICV_4 $T=413120 270880 0 0 $X=412830 $Y=270645
X689 1 2 ICV_4 $T=434400 247360 0 0 $X=434110 $Y=247125
X690 1 2 ICV_4 $T=455120 239520 1 0 $X=454830 $Y=235310
X691 268 264 257 2 1 1071 DFCNQD1BWP7T $T=197520 231680 1 180 $X=184910 $Y=231445
X692 268 1106 257 2 1 1084 DFCNQD1BWP7T $T=218240 239520 1 180 $X=205630 $Y=239285
X693 268 1107 257 2 1 1103 DFCNQD1BWP7T $T=218240 255200 0 180 $X=205630 $Y=250990
X694 268 1108 287 2 1 1067 DFCNQD1BWP7T $T=218240 263040 0 180 $X=205630 $Y=258830
X695 268 289 257 2 1 1100 DFCNQD1BWP7T $T=218800 231680 1 180 $X=206190 $Y=231445
X696 268 1111 287 2 1 1101 DFCNQD1BWP7T $T=220480 263040 1 180 $X=207870 $Y=262805
X697 268 1112 287 2 1 1038 DFCNQD1BWP7T $T=220480 270880 0 180 $X=207870 $Y=266670
X698 268 1116 287 2 1 1065 DFCNQD1BWP7T $T=224960 286560 0 180 $X=212350 $Y=282350
X699 268 297 257 2 1 1088 DFCNQD1BWP7T $T=226640 239520 0 180 $X=214030 $Y=235310
X700 268 298 287 2 1 1105 DFCNQD1BWP7T $T=227200 270880 1 180 $X=214590 $Y=270645
X701 268 1123 287 2 1 1083 DFCNQD1BWP7T $T=231120 294400 0 180 $X=218510 $Y=290190
X702 268 1124 287 2 1 1109 DFCNQD1BWP7T $T=234480 270880 0 180 $X=221870 $Y=266670
X703 268 1154 287 2 1 1138 DFCNQD1BWP7T $T=260800 270880 1 180 $X=248190 $Y=270645
X704 268 1183 417 2 1 1157 DFCNQD1BWP7T $T=290480 294400 1 0 $X=290190 $Y=290190
X705 268 1187 417 2 1 425 DFCNQD1BWP7T $T=294960 286560 0 0 $X=294670 $Y=286325
X706 468 1268 282 2 1 1266 DFCNQD1BWP7T $T=445040 263040 0 180 $X=432430 $Y=258830
X707 468 1273 282 2 1 1267 DFCNQD1BWP7T $T=448960 255200 1 180 $X=436350 $Y=254965
X973 1 2 ICV_8 $T=20000 263040 0 0 $X=19710 $Y=262805
X974 1 2 ICV_8 $T=20000 278720 1 0 $X=19710 $Y=274510
X975 1 2 ICV_8 $T=34000 255200 1 0 $X=33710 $Y=250990
X976 1 2 ICV_8 $T=34000 278720 0 0 $X=33710 $Y=278485
X977 1 2 ICV_8 $T=76000 270880 0 0 $X=75710 $Y=270645
X978 1 2 ICV_8 $T=118000 247360 0 0 $X=117710 $Y=247125
X979 1 2 ICV_8 $T=118000 263040 0 0 $X=117710 $Y=262805
X980 1 2 ICV_8 $T=118000 270880 0 0 $X=117710 $Y=270645
X981 1 2 ICV_8 $T=118000 278720 1 0 $X=117710 $Y=274510
X982 1 2 ICV_8 $T=160000 231680 0 0 $X=159710 $Y=231445
X983 1 2 ICV_8 $T=160000 239520 1 0 $X=159710 $Y=235310
X984 1 2 ICV_8 $T=160000 239520 0 0 $X=159710 $Y=239285
X985 1 2 ICV_8 $T=160000 255200 1 0 $X=159710 $Y=250990
X986 1 2 ICV_8 $T=160000 255200 0 0 $X=159710 $Y=254965
X987 1 2 ICV_8 $T=160000 263040 1 0 $X=159710 $Y=258830
X988 1 2 ICV_8 $T=160000 263040 0 0 $X=159710 $Y=262805
X989 1 2 ICV_8 $T=160000 270880 1 0 $X=159710 $Y=266670
X990 1 2 ICV_8 $T=160000 278720 0 0 $X=159710 $Y=278485
X991 1 2 ICV_8 $T=160000 286560 0 0 $X=159710 $Y=286325
X992 1 2 ICV_8 $T=160000 294400 1 0 $X=159710 $Y=290190
X993 1 2 ICV_8 $T=202000 239520 0 0 $X=201710 $Y=239285
X994 1 2 ICV_8 $T=202000 255200 1 0 $X=201710 $Y=250990
X995 1 2 ICV_8 $T=202000 263040 1 0 $X=201710 $Y=258830
X996 1 2 ICV_8 $T=244000 247360 1 0 $X=243710 $Y=243150
X997 1 2 ICV_8 $T=286000 263040 0 0 $X=285710 $Y=262805
X998 1 2 ICV_8 $T=286000 270880 1 0 $X=285710 $Y=266670
X999 1 2 ICV_8 $T=286000 278720 0 0 $X=285710 $Y=278485
X1000 1 2 ICV_8 $T=328000 255200 0 0 $X=327710 $Y=254965
X1001 1 2 ICV_8 $T=328000 278720 0 0 $X=327710 $Y=278485
X1002 1 2 ICV_8 $T=370000 231680 0 0 $X=369710 $Y=231445
X1003 1 2 ICV_8 $T=370000 255200 1 0 $X=369710 $Y=250990
X1004 1 2 ICV_8 $T=412000 239520 0 0 $X=411710 $Y=239285
X1005 1 2 ICV_8 $T=454000 231680 0 0 $X=453710 $Y=231445
X1006 1 2 ICV_8 $T=454000 263040 1 0 $X=453710 $Y=258830
X1007 1 2 ICV_9 $T=20000 231680 0 0 $X=19710 $Y=231445
X1008 1 2 ICV_9 $T=20000 270880 1 0 $X=19710 $Y=266670
X1009 1 2 ICV_9 $T=20000 294400 1 0 $X=19710 $Y=290190
X1010 1 2 ICV_9 $T=34000 231680 0 0 $X=33710 $Y=231445
X1011 1 2 ICV_9 $T=34000 263040 0 0 $X=33710 $Y=262805
X1012 1 2 ICV_9 $T=34000 270880 1 0 $X=33710 $Y=266670
X1013 1 2 ICV_9 $T=34000 270880 0 0 $X=33710 $Y=270645
X1014 1 2 ICV_9 $T=34000 278720 1 0 $X=33710 $Y=274510
X1015 1 2 ICV_9 $T=118000 278720 0 0 $X=117710 $Y=278485
X1016 1 2 ICV_9 $T=118000 294400 1 0 $X=117710 $Y=290190
X1017 1 2 ICV_9 $T=160000 247360 0 0 $X=159710 $Y=247125
X1018 1 2 ICV_9 $T=202000 247360 1 0 $X=201710 $Y=243150
X1019 1 2 ICV_9 $T=202000 247360 0 0 $X=201710 $Y=247125
X1020 1 2 ICV_9 $T=202000 255200 0 0 $X=201710 $Y=254965
X1021 1 2 ICV_9 $T=202000 263040 0 0 $X=201710 $Y=262805
X1022 1 2 ICV_9 $T=202000 270880 1 0 $X=201710 $Y=266670
X1023 1 2 ICV_9 $T=202000 278720 1 0 $X=201710 $Y=274510
X1024 1 2 ICV_9 $T=202000 286560 0 0 $X=201710 $Y=286325
X1025 1 2 ICV_9 $T=244000 255200 1 0 $X=243710 $Y=250990
X1026 1 2 ICV_9 $T=244000 286560 1 0 $X=243710 $Y=282350
X1027 1 2 ICV_9 $T=244000 286560 0 0 $X=243710 $Y=286325
X1028 1 2 ICV_9 $T=286000 247360 0 0 $X=285710 $Y=247125
X1029 1 2 ICV_9 $T=286000 255200 1 0 $X=285710 $Y=250990
X1030 1 2 ICV_9 $T=286000 255200 0 0 $X=285710 $Y=254965
X1031 1 2 ICV_9 $T=286000 270880 0 0 $X=285710 $Y=270645
X1032 1 2 ICV_9 $T=286000 286560 1 0 $X=285710 $Y=282350
X1033 1 2 ICV_9 $T=328000 239520 0 0 $X=327710 $Y=239285
X1034 1 2 ICV_9 $T=328000 263040 1 0 $X=327710 $Y=258830
X1035 1 2 ICV_9 $T=328000 286560 1 0 $X=327710 $Y=282350
X1036 1 2 ICV_9 $T=370000 239520 0 0 $X=369710 $Y=239285
X1037 1 2 ICV_9 $T=370000 247360 1 0 $X=369710 $Y=243150
X1038 1 2 ICV_9 $T=370000 255200 0 0 $X=369710 $Y=254965
X1039 1 2 ICV_9 $T=370000 263040 0 0 $X=369710 $Y=262805
X1040 1 2 ICV_9 $T=370000 270880 0 0 $X=369710 $Y=270645
X1041 1 2 ICV_9 $T=370000 278720 0 0 $X=369710 $Y=278485
X1042 1 2 ICV_9 $T=412000 239520 1 0 $X=411710 $Y=235310
X1043 1 2 ICV_9 $T=412000 263040 0 0 $X=411710 $Y=262805
X1044 1 2 ICV_9 $T=454000 247360 1 0 $X=453710 $Y=243150
X1045 1 2 ICV_9 $T=454000 263040 0 0 $X=453710 $Y=262805
X1046 1 2 ICV_9 $T=454000 278720 0 0 $X=453710 $Y=278485
X1047 1 2 ICV_9 $T=454000 286560 1 0 $X=453710 $Y=282350
X1048 1 2 ICV_9 $T=454000 286560 0 0 $X=453710 $Y=286325
X1049 1 2 ICV_9 $T=454000 294400 1 0 $X=453710 $Y=290190
X1092 1 2 ICV_13 $T=30640 247360 0 0 $X=30350 $Y=247125
X1093 1 2 ICV_13 $T=35120 239520 0 0 $X=34830 $Y=239285
X1094 1 2 ICV_13 $T=53600 286560 1 0 $X=53310 $Y=282350
X1095 1 2 ICV_13 $T=54720 255200 1 0 $X=54430 $Y=250990
X1096 1 2 ICV_13 $T=63120 270880 1 0 $X=62830 $Y=266670
X1097 1 2 ICV_13 $T=67040 278720 0 0 $X=66750 $Y=278485
X1098 1 2 ICV_13 $T=72640 255200 0 0 $X=72350 $Y=254965
X1099 1 2 ICV_13 $T=77120 239520 1 0 $X=76830 $Y=235310
X1100 1 2 ICV_13 $T=96720 286560 1 0 $X=96430 $Y=282350
X1101 1 2 ICV_13 $T=135360 278720 1 0 $X=135070 $Y=274510
X1102 1 2 ICV_13 $T=139840 239520 0 0 $X=139550 $Y=239285
X1103 1 2 ICV_13 $T=142640 247360 0 0 $X=142350 $Y=247125
X1104 1 2 ICV_13 $T=156640 247360 0 0 $X=156350 $Y=247125
X1105 1 2 ICV_13 $T=171760 255200 1 0 $X=171470 $Y=250990
X1106 1 2 ICV_13 $T=179040 270880 0 0 $X=178750 $Y=270645
X1107 1 2 ICV_13 $T=181840 231680 0 0 $X=181550 $Y=231445
X1108 1 2 ICV_13 $T=198640 239520 0 0 $X=198350 $Y=239285
X1109 1 2 ICV_13 $T=203120 294400 1 0 $X=202830 $Y=290190
X1110 1 2 ICV_13 $T=207600 255200 0 0 $X=207310 $Y=254965
X1111 1 2 ICV_13 $T=207600 278720 1 0 $X=207310 $Y=274510
X1112 1 2 ICV_13 $T=217680 278720 1 0 $X=217390 $Y=274510
X1113 1 2 ICV_13 $T=240640 231680 0 0 $X=240350 $Y=231445
X1114 1 2 ICV_13 $T=240640 263040 0 0 $X=240350 $Y=262805
X1115 1 2 ICV_13 $T=240640 278720 0 0 $X=240350 $Y=278485
X1116 1 2 ICV_13 $T=249600 286560 1 0 $X=249310 $Y=282350
X1117 1 2 ICV_13 $T=272000 255200 1 0 $X=271710 $Y=250990
X1118 1 2 ICV_13 $T=282640 239520 1 0 $X=282350 $Y=235310
X1119 1 2 ICV_13 $T=282640 278720 1 0 $X=282350 $Y=274510
X1120 1 2 ICV_13 $T=292160 270880 1 0 $X=291870 $Y=266670
X1121 1 2 ICV_13 $T=294960 255200 0 0 $X=294670 $Y=254965
X1122 1 2 ICV_13 $T=311760 294400 1 0 $X=311470 $Y=290190
X1123 1 2 ICV_13 $T=319600 270880 0 0 $X=319310 $Y=270645
X1124 1 2 ICV_13 $T=329120 247360 0 0 $X=328830 $Y=247125
X1125 1 2 ICV_13 $T=385120 294400 1 0 $X=384830 $Y=290190
X1126 1 2 ICV_13 $T=417600 263040 0 0 $X=417310 $Y=262805
X1127 1 2 ICV_13 $T=424320 239520 0 0 $X=424030 $Y=239285
X1128 1 2 ICV_13 $T=450640 231680 0 0 $X=450350 $Y=231445
X1129 1 2 ICV_13 $T=450640 278720 0 0 $X=450350 $Y=278485
X1130 1 2 ICV_13 $T=450640 286560 1 0 $X=450350 $Y=282350
X1131 1 2 ICV_13 $T=450640 286560 0 0 $X=450350 $Y=286325
X1132 1 2 ICV_13 $T=455120 247360 0 0 $X=454830 $Y=247125
X1133 1 2 ICV_13 $T=455120 270880 1 0 $X=454830 $Y=266670
X1134 1 2 ICV_13 $T=459600 263040 0 0 $X=459310 $Y=262805
X1135 225 1050 2 1050 1053 225 1 MAOI22D1BWP7T $T=179040 270880 1 180 $X=174270 $Y=270645
X1136 1024 226 2 226 1074 1024 1 MAOI22D1BWP7T $T=177920 263040 0 0 $X=177630 $Y=262805
X1137 1181 1186 2 1186 1185 1181 1 MAOI22D1BWP7T $T=298320 247360 0 180 $X=293550 $Y=243150
X1138 447 445 2 447 446 445 1 MAOI22D1BWP7T $T=317920 239520 0 180 $X=313150 $Y=235310
X1139 1201 449 2 449 1188 1201 1 MAOI22D1BWP7T $T=319040 255200 1 180 $X=314270 $Y=254965
X1140 473 477 2 477 1207 473 1 MAOI22D1BWP7T $T=333040 239520 1 0 $X=332750 $Y=235310
X1141 1214 523 2 523 1232 1214 1 MAOI22D1BWP7T $T=374480 270880 1 0 $X=374190 $Y=266670
X1142 589 587 2 589 1263 587 1 MAOI22D1BWP7T $T=426000 263040 1 180 $X=421230 $Y=262805
X1143 1184 274 1 1106 407 2 IOA21D0BWP7T $T=294400 239520 1 180 $X=290750 $Y=239285
X1144 8 1 2 862 INVD1BWP7T $T=31200 286560 0 180 $X=29230 $Y=282350
X1145 29 1 2 872 INVD1BWP7T $T=40160 278720 1 0 $X=39870 $Y=274510
X1146 892 1 2 893 INVD1BWP7T $T=51360 247360 1 0 $X=51070 $Y=243150
X1147 860 1 2 889 INVD1BWP7T $T=53040 255200 1 0 $X=52750 $Y=250990
X1148 878 1 2 55 INVD1BWP7T $T=53600 239520 1 0 $X=53310 $Y=235310
X1149 867 1 2 59 INVD1BWP7T $T=56960 270880 0 0 $X=56670 $Y=270645
X1150 910 1 2 909 INVD1BWP7T $T=63680 263040 0 0 $X=63390 $Y=262805
X1151 863 1 2 929 INVD1BWP7T $T=66480 270880 1 0 $X=66190 $Y=266670
X1152 902 1 2 891 INVD1BWP7T $T=73200 255200 0 180 $X=71230 $Y=250990
X1153 4 1 2 907 INVD1BWP7T $T=80480 255200 0 0 $X=80190 $Y=254965
X1154 969 1 2 882 INVD1BWP7T $T=98400 247360 1 180 $X=96430 $Y=247125
X1155 933 1 2 967 INVD1BWP7T $T=108480 255200 1 0 $X=108190 $Y=250990
X1156 106 1 2 997 INVD1BWP7T $T=121920 263040 0 0 $X=121630 $Y=262805
X1157 1007 1 2 144 INVD1BWP7T $T=133680 270880 0 180 $X=131710 $Y=266670
X1158 171 1 2 1002 INVD1BWP7T $T=137600 255200 0 0 $X=137310 $Y=254965
X1159 155 1 2 1001 INVD1BWP7T $T=147680 247360 1 180 $X=145710 $Y=247125
X1160 192 1 2 1040 INVD1BWP7T $T=154400 286560 0 0 $X=154110 $Y=286325
X1161 225 1 2 223 INVD1BWP7T $T=181280 278720 1 0 $X=180990 $Y=274510
X1162 239 1 2 1068 INVD1BWP7T $T=185760 247360 1 180 $X=183790 $Y=247125
X1163 1089 1 2 1080 INVD1BWP7T $T=189680 270880 1 180 $X=187710 $Y=270645
X1164 348 1 2 342 INVD1BWP7T $T=255200 278720 0 180 $X=253230 $Y=274510
X1165 273 1 2 368 INVD1BWP7T $T=268640 286560 1 0 $X=268350 $Y=282350
X1166 456 1 2 474 INVD1BWP7T $T=334720 270880 0 180 $X=332750 $Y=266670
X1167 563 1 2 566 INVD1BWP7T $T=400800 255200 1 0 $X=400510 $Y=250990
X1168 1 2 ICV_14 $T=28400 247360 1 0 $X=28110 $Y=243150
X1169 1 2 ICV_14 $T=46320 239520 0 0 $X=46030 $Y=239285
X1170 1 2 ICV_14 $T=47440 255200 0 0 $X=47150 $Y=254965
X1171 1 2 ICV_14 $T=106800 247360 1 0 $X=106510 $Y=243150
X1172 1 2 ICV_14 $T=129200 255200 0 0 $X=128910 $Y=254965
X1173 1 2 ICV_14 $T=154400 255200 1 0 $X=154110 $Y=250990
X1174 1 2 ICV_14 $T=218240 255200 1 0 $X=217950 $Y=250990
X1175 1 2 ICV_14 $T=263600 286560 0 0 $X=263310 $Y=286325
X1176 1 2 ICV_14 $T=269760 270880 1 0 $X=269470 $Y=266670
X1177 1 2 ICV_14 $T=271440 286560 0 0 $X=271150 $Y=286325
X1178 1 2 ICV_14 $T=299440 247360 0 0 $X=299150 $Y=247125
X1179 1 2 ICV_14 $T=308960 239520 0 0 $X=308670 $Y=239285
X1180 1 2 ICV_14 $T=322400 270880 1 0 $X=322110 $Y=266670
X1181 1 2 ICV_14 $T=356000 239520 1 0 $X=355710 $Y=235310
X1182 1 2 ICV_14 $T=371120 286560 1 0 $X=370830 $Y=282350
X1183 1 2 ICV_14 $T=406400 263040 0 0 $X=406110 $Y=262805
X1184 1 2 ICV_14 $T=406400 294400 1 0 $X=406110 $Y=290190
X1185 1 2 ICV_14 $T=435520 231680 0 0 $X=435230 $Y=231445
X1186 1 2 ICV_14 $T=435520 263040 0 0 $X=435230 $Y=262805
X1187 1 2 ICV_14 $T=448400 239520 0 0 $X=448110 $Y=239285
X1188 1 2 ICV_14 $T=462400 286560 0 0 $X=462110 $Y=286325
X1189 503 381 1 2 BUFFD10BWP7T $T=356000 278720 0 180 $X=345070 $Y=274510
X1190 1109 281 1 2 BUFFD2BWP7T $T=212080 247360 1 180 $X=208430 $Y=247125
X1191 457 436 1 2 BUFFD2BWP7T $T=318480 294400 0 180 $X=314830 $Y=290190
X1192 638 639 1 2 BUFFD2BWP7T $T=447280 286560 0 0 $X=446990 $Y=286325
X1193 678 661 1 2 BUFFD2BWP7T $T=470800 270880 0 180 $X=467150 $Y=266670
X1194 1 2 DCAP16BWP7T $T=119120 239520 1 0 $X=118830 $Y=235310
X1195 1 2 DCAP16BWP7T $T=119120 247360 1 0 $X=118830 $Y=243150
X1196 1 2 DCAP16BWP7T $T=148800 263040 0 0 $X=148510 $Y=262805
X1197 1 2 DCAP16BWP7T $T=191360 263040 1 0 $X=191070 $Y=258830
X1198 1 2 DCAP16BWP7T $T=218800 231680 0 0 $X=218510 $Y=231445
X1199 1 2 DCAP16BWP7T $T=231680 263040 0 0 $X=231390 $Y=262805
X1200 1 2 DCAP16BWP7T $T=262480 255200 0 0 $X=262190 $Y=254965
X1201 1 2 DCAP16BWP7T $T=302800 294400 1 0 $X=302510 $Y=290190
X1202 1 2 DCAP16BWP7T $T=317920 239520 1 0 $X=317630 $Y=235310
X1203 1 2 DCAP16BWP7T $T=318480 294400 1 0 $X=318190 $Y=290190
X1204 1 2 DCAP16BWP7T $T=319040 255200 0 0 $X=318750 $Y=254965
X1205 1 2 DCAP16BWP7T $T=329120 270880 0 0 $X=328830 $Y=270645
X1206 1 2 DCAP16BWP7T $T=352080 255200 1 0 $X=351790 $Y=250990
X1207 1 2 DCAP16BWP7T $T=356000 278720 1 0 $X=355710 $Y=274510
X1208 1 2 DCAP16BWP7T $T=359920 247360 1 0 $X=359630 $Y=243150
X1209 1 2 DCAP16BWP7T $T=359920 270880 0 0 $X=359630 $Y=270645
X1210 1 2 DCAP16BWP7T $T=371120 263040 1 0 $X=370830 $Y=258830
X1211 1 2 DCAP16BWP7T $T=385680 263040 0 0 $X=385390 $Y=262805
X1212 1 2 DCAP16BWP7T $T=401360 247360 0 0 $X=401070 $Y=247125
X1213 1 2 DCAP16BWP7T $T=401360 278720 0 0 $X=401070 $Y=278485
X1214 1 2 DCAP16BWP7T $T=413120 247360 1 0 $X=412830 $Y=243150
X1215 1 2 DCAP16BWP7T $T=413120 278720 0 0 $X=412830 $Y=278485
X1216 1 2 DCAP16BWP7T $T=425440 247360 0 0 $X=425150 $Y=247125
X1217 1 2 DCAP16BWP7T $T=425440 286560 1 0 $X=425150 $Y=282350
X1218 1 2 DCAP16BWP7T $T=441680 278720 0 0 $X=441390 $Y=278485
X1219 1 2 DCAP16BWP7T $T=441680 286560 1 0 $X=441390 $Y=282350
X1220 1 2 DCAP16BWP7T $T=443360 247360 1 0 $X=443070 $Y=243150
X1221 1 2 DCAP16BWP7T $T=444480 247360 0 0 $X=444190 $Y=247125
X1222 1 2 DCAP16BWP7T $T=444480 270880 1 0 $X=444190 $Y=266670
X1223 1 2 DCAP16BWP7T $T=445040 263040 1 0 $X=444750 $Y=258830
X1224 5 1 2 861 CKND1BWP7T $T=25600 286560 1 0 $X=25310 $Y=282350
X1225 921 1 2 931 CKND1BWP7T $T=88880 247360 1 180 $X=86910 $Y=247125
X1226 211 1 2 1045 CKND1BWP7T $T=163920 294400 1 0 $X=163630 $Y=290190
X1227 216 1 2 1044 CKND1BWP7T $T=166720 270880 1 180 $X=164750 $Y=270645
X1228 246 1 2 1075 CKND1BWP7T $T=184640 278720 0 180 $X=182670 $Y=274510
X1229 608 1 2 612 CKND1BWP7T $T=433840 231680 0 0 $X=433550 $Y=231445
X1230 1267 1 2 310 BUFFD3BWP7T $T=439440 247360 1 0 $X=439150 $Y=243150
X1231 671 447 1 2 BUFFD12BWP7T $T=470800 255200 0 180 $X=458190 $Y=250990
X1232 1110 283 277 1 2 CKXOR2D4BWP7T $T=218800 294400 0 180 $X=206190 $Y=290190
X1233 562 1245 545 1 2 CKXOR2D4BWP7T $T=401360 247360 1 180 $X=388750 $Y=247125
X1234 620 611 892 1 2 CKXOR2D4BWP7T $T=441680 278720 1 180 $X=429070 $Y=278485
X1235 168 1013 2 944 1 163 1029 AOI22D1BWP7T $T=138720 286560 1 0 $X=138430 $Y=282350
X1236 192 198 2 1040 1 197 1023 AOI22D1BWP7T $T=157200 278720 0 180 $X=152990 $Y=274510
X1237 1039 198 2 1034 1 197 1042 AOI22D1BWP7T $T=153280 286560 1 0 $X=152990 $Y=282350
X1238 208 1040 2 201 1 192 193 AOI22D1BWP7T $T=157200 294400 0 180 $X=152990 $Y=290190
X1239 1044 212 2 216 1 217 1051 AOI22D1BWP7T $T=163920 270880 1 0 $X=163630 $Y=266670
X1240 1045 212 2 211 1 217 1054 AOI22D1BWP7T $T=163920 278720 0 0 $X=163630 $Y=278485
X1241 1048 1043 2 210 1 1049 1052 AOI22D1BWP7T $T=165600 239520 0 0 $X=165310 $Y=239285
X1242 225 239 2 223 1 1068 1046 AOI22D1BWP7T $T=179600 255200 0 180 $X=175390 $Y=250990
X1243 198 1056 2 197 1 213 1073 AOI22D1BWP7T $T=177360 278720 1 0 $X=177070 $Y=274510
X1244 225 1075 2 223 1 246 243 AOI22D1BWP7T $T=180160 278720 0 0 $X=179870 $Y=278485
X1245 1081 1075 2 1061 1 246 1079 AOI22D1BWP7T $T=186320 270880 1 180 $X=182110 $Y=270645
X1246 309 292 2 1113 1 312 1131 AOI22D1BWP7T $T=228880 239520 0 0 $X=228590 $Y=239285
X1247 1130 331 2 313 1 316 1140 AOI22D1BWP7T $T=247920 247360 1 0 $X=247630 $Y=243150
X1248 1139 331 2 330 1 316 1137 AOI22D1BWP7T $T=252400 231680 1 180 $X=248190 $Y=231445
X1249 340 1153 2 349 1 1136 353 AOI22D1BWP7T $T=259680 270880 0 180 $X=255470 $Y=266670
X1250 360 273 2 1143 1 368 382 AOI22D1BWP7T $T=264160 278720 0 0 $X=263870 $Y=278485
X1251 381 396 2 391 1 389 1174 AOI22D1BWP7T $T=280400 231680 1 180 $X=276190 $Y=231445
X1252 1223 502 2 1222 1 500 488 AOI22D1BWP7T $T=356000 239520 0 180 $X=351790 $Y=235310
X1253 1249 563 2 1250 1 566 1252 AOI22D1BWP7T $T=398560 263040 1 0 $X=398270 $Y=258830
X1254 1251 563 2 569 1 566 1255 AOI22D1BWP7T $T=402480 263040 0 0 $X=402190 $Y=262805
X1255 381 575 2 450 1 572 573 AOI22D1BWP7T $T=408080 270880 1 180 $X=403870 $Y=270645
X1256 448 615 2 450 1 610 607 AOI22D1BWP7T $T=437760 286560 1 180 $X=433550 $Y=286325
X1257 448 565 2 450 1 627 636 AOI22D1BWP7T $T=442240 270880 0 0 $X=441950 $Y=270645
X1258 25 16 2 872 28 1 OAI21D1BWP7T $T=37920 278720 0 0 $X=37630 $Y=278485
X1259 344 1140 2 1142 1148 1 OAI21D1BWP7T $T=254640 255200 1 180 $X=250990 $Y=254965
X1260 323 1167 2 362 1164 1 OAI21D1BWP7T $T=261360 255200 1 0 $X=261070 $Y=250990
X1261 376 1173 2 1174 378 1 OAI21D1BWP7T $T=270320 247360 0 0 $X=270030 $Y=247125
X1262 376 1178 2 406 1111 1 OAI21D1BWP7T $T=278160 247360 0 0 $X=277870 $Y=247125
X1263 409 1175 2 1182 414 1 OAI21D1BWP7T $T=292160 278720 1 0 $X=291870 $Y=274510
X1264 323 1202 2 452 1191 1 OAI21D1BWP7T $T=314560 239520 0 0 $X=314270 $Y=239285
X1265 443 451 1 2 BUFFD8BWP7T $T=311760 231680 0 0 $X=311470 $Y=231445
X1266 282 257 1 2 BUFFD6BWP7T $T=210960 255200 0 0 $X=210670 $Y=254965
X1267 851 847 2 1 INVD2BWP7T $T=23360 263040 0 180 $X=20830 $Y=258830
X1268 856 25 2 1 INVD2BWP7T $T=39040 263040 1 0 $X=38750 $Y=258830
X1269 37 20 2 1 INVD2BWP7T $T=46320 239520 1 180 $X=43790 $Y=239285
X1270 65 879 2 1 INVD2BWP7T $T=67040 286560 0 180 $X=64510 $Y=282350
X1271 846 916 2 1 INVD2BWP7T $T=111280 239520 0 0 $X=110990 $Y=239285
X1272 985 110 2 1 INVD2BWP7T $T=125840 263040 1 180 $X=123310 $Y=262805
X1273 915 908 2 1 INVD2BWP7T $T=133680 255200 0 180 $X=131150 $Y=250990
X1274 963 868 2 1 INVD2BWP7T $T=134800 247360 0 180 $X=132270 $Y=243150
X1275 309 347 2 1 INVD2BWP7T $T=253520 286560 1 0 $X=253230 $Y=282350
X1276 1157 383 2 1 INVD2BWP7T $T=272560 263040 1 0 $X=272270 $Y=258830
X1277 393 384 2 1 INVD2BWP7T $T=278160 247360 0 180 $X=275630 $Y=243150
X1278 387 513 2 1 INVD2BWP7T $T=364960 286560 0 180 $X=362430 $Y=282350
X1279 541 543 2 1 INVD2BWP7T $T=387360 270880 1 0 $X=387070 $Y=266670
X1280 603 557 2 1 INVD2BWP7T $T=429920 239520 1 180 $X=427390 $Y=239285
X1281 615 574 2 1 INVD2BWP7T $T=439440 294400 0 180 $X=436910 $Y=290190
X1282 611 578 2 1 INVD2BWP7T $T=446720 294400 0 180 $X=444190 $Y=290190
X1283 199 242 1 2 1077 CKXOR2D1BWP7T $T=177360 286560 0 0 $X=177070 $Y=286325
X1284 213 241 1 2 1072 CKXOR2D1BWP7T $T=184080 247360 1 180 $X=178750 $Y=247125
X1285 223 238 1 2 1049 CKXOR2D1BWP7T $T=184640 247360 0 180 $X=179310 $Y=243150
X1286 206 247 1 2 1050 CKXOR2D1BWP7T $T=181280 270880 1 0 $X=180990 $Y=266670
X1287 1050 1080 1 2 1066 CKXOR2D1BWP7T $T=191360 263040 0 180 $X=186030 $Y=258830
X1288 1049 1091 1 2 269 CKXOR2D1BWP7T $T=210960 270880 1 180 $X=205630 $Y=270645
X1289 290 292 1 2 1113 CKXOR2D1BWP7T $T=216560 247360 0 0 $X=216270 $Y=247125
X1290 293 292 1 2 303 CKXOR2D1BWP7T $T=219920 239520 0 0 $X=219630 $Y=239285
X1291 1127 321 1 2 1134 CKXOR2D1BWP7T $T=234480 270880 0 0 $X=234190 $Y=270645
X1292 1117 327 1 2 1136 CKXOR2D1BWP7T $T=236160 263040 1 0 $X=235870 $Y=258830
X1293 368 300 1 2 422 CKXOR2D1BWP7T $T=292160 286560 1 0 $X=291870 $Y=282350
X1294 435 1199 1 2 1195 CKXOR2D1BWP7T $T=305040 247360 0 0 $X=304750 $Y=247125
X1295 1195 444 1 2 1196 CKXOR2D1BWP7T $T=308960 270880 1 0 $X=308670 $Y=266670
X1296 499 366 1 2 495 CKXOR2D1BWP7T $T=351520 286560 0 180 $X=346190 $Y=282350
X1297 1237 547 1 2 1235 CKXOR2D1BWP7T $T=392960 255200 0 180 $X=387630 $Y=250990
X1298 1047 1036 224 1 2 CKXOR2D2BWP7T $T=163920 263040 1 0 $X=163630 $Y=258830
X1299 1072 1063 248 1 2 CKXOR2D2BWP7T $T=179040 239520 1 0 $X=178750 $Y=235310
X1300 1049 1090 272 1 2 CKXOR2D2BWP7T $T=193040 270880 0 0 $X=192750 $Y=270645
X1301 288 280 278 1 2 CKXOR2D2BWP7T $T=214320 286560 1 180 $X=207870 $Y=286325
X1302 310 1121 299 1 2 CKXOR2D2BWP7T $T=231120 247360 0 180 $X=224670 $Y=243150
X1303 1164 1157 350 1 2 CKXOR2D2BWP7T $T=263600 286560 1 180 $X=257150 $Y=286325
X1304 1191 425 420 1 2 CKXOR2D2BWP7T $T=303920 255200 0 180 $X=297470 $Y=250990
X1305 441 436 432 1 2 CKXOR2D2BWP7T $T=310640 286560 0 180 $X=304190 $Y=282350
X1306 2 1 DCAP32BWP7T $T=292160 263040 0 0 $X=291870 $Y=262805
X1307 2 1 DCAP32BWP7T $T=349840 231680 0 0 $X=349550 $Y=231445
X1308 1052 1084 259 1078 262 1 2 XNR4D1BWP7T $T=184640 247360 1 0 $X=184350 $Y=243150
X1309 279 1 2 387 BUFFD5BWP7T $T=272560 239520 0 0 $X=272270 $Y=239285
X1310 1141 1145 338 340 1 2 OAI21D0BWP7T $T=251280 239520 0 0 $X=250990 $Y=239285
X1311 1158 1165 1162 340 1 2 OAI21D0BWP7T $T=263600 247360 1 0 $X=263310 $Y=243150
X1312 351 1163 375 1170 1 2 OAI21D0BWP7T $T=266960 247360 1 0 $X=266670 $Y=243150
X1313 430 1197 433 427 1 2 OAI21D0BWP7T $T=307840 247360 1 0 $X=307550 $Y=243150
X1314 1216 1217 497 427 1 2 OAI21D0BWP7T $T=348720 239520 0 0 $X=348430 $Y=239285
X1315 521 538 532 1238 1 2 OAI21D0BWP7T $T=383440 239520 0 180 $X=380350 $Y=235310
X1316 1255 1259 580 427 1 2 OAI21D0BWP7T $T=416480 247360 0 0 $X=416190 $Y=247125
X1317 1256 1254 582 1262 1 2 OAI21D0BWP7T $T=421520 239520 0 0 $X=421230 $Y=239285
X1318 1261 1264 591 340 1 2 OAI21D0BWP7T $T=422640 286560 1 0 $X=422350 $Y=282350
X1319 180 185 1035 1033 204 1 2 XNR4D0BWP7T $T=144320 247360 1 0 $X=144030 $Y=243150
X1320 1023 1026 1036 1038 1041 1 2 XNR4D0BWP7T $T=144320 263040 1 0 $X=144030 $Y=258830
X1321 1024 1027 1037 193 205 1 2 XNR4D0BWP7T $T=144320 270880 1 0 $X=144030 $Y=266670
X1322 1067 230 1055 220 210 1 2 XNR4D0BWP7T $T=176800 263040 1 180 $X=163630 $Y=262805
X1323 215 1054 1063 1033 238 1 2 XNR4D0BWP7T $T=165600 239520 1 0 $X=165310 $Y=235310
X1324 1070 1064 1058 1051 1050 1 2 XNR4D0BWP7T $T=179040 247360 1 180 $X=165870 $Y=247125
X1325 1053 227 234 1042 241 1 2 XNR4D0BWP7T $T=167280 294400 1 0 $X=166990 $Y=290190
X1326 1076 251 1090 255 262 1 2 XNR4D0BWP7T $T=181280 294400 1 0 $X=180990 $Y=290190
X1327 1103 1074 1093 216 1080 1 2 XNR4D0BWP7T $T=199200 255200 1 180 $X=186030 $Y=254965
X1328 1101 1073 1094 205 1050 1 2 XNR4D0BWP7T $T=199200 270880 0 180 $X=186030 $Y=266670
X1329 1035 1027 231 1051 237 1 2 XNR4D2BWP7T $T=164480 247360 1 0 $X=164190 $Y=243150
X1330 221 1041 235 1042 242 1 2 XNR4D2BWP7T $T=167280 286560 1 0 $X=166990 $Y=282350
X1331 222 1060 236 1024 1050 1 2 XNR4D2BWP7T $T=167840 270880 1 0 $X=167550 $Y=266670
X1332 1057 1071 232 1060 226 1 2 XNR4D2BWP7T $T=182960 239520 1 180 $X=169230 $Y=239285
X1333 1055 1046 240 1066 241 1 2 XNR4D2BWP7T $T=170080 263040 1 0 $X=169790 $Y=258830
X1334 228 1066 244 1072 1068 1 2 XNR4D2BWP7T $T=172320 255200 0 0 $X=172030 $Y=254965
X1335 1076 250 256 1069 1061 1 2 XNR4D2BWP7T $T=181280 286560 1 0 $X=180990 $Y=282350
X1336 211 1083 260 1077 269 1 2 XNR4D2BWP7T $T=184080 286560 0 0 $X=183790 $Y=286325
X1337 1057 1085 261 1073 258 1 2 XNR4D2BWP7T $T=184640 255200 1 0 $X=184350 $Y=250990
X1338 239 1088 263 266 1074 1 2 XNR4D2BWP7T $T=185200 239520 0 0 $X=184910 $Y=239285
X1339 1079 253 265 1078 1069 1 2 XNR4D2BWP7T $T=185760 247360 0 0 $X=185470 $Y=247125
X1340 1087 267 1092 1034 1080 1 2 XNR4D2BWP7T $T=199200 278720 0 180 $X=185470 $Y=274510
X1341 270 1105 286 1077 247 1 2 XNR4D2BWP7T $T=220480 278720 1 180 $X=206750 $Y=278485
X1342 213 1026 1056 1 2 1061 MUX2ND1BWP7T $T=166160 255200 0 0 $X=165870 $Y=254965
X1343 1171 1135 1168 1 2 1166 MUX2ND1BWP7T $T=271440 263040 0 180 $X=264990 $Y=258830
X1344 484 480 1214 1 2 1212 MUX2ND1BWP7T $T=336400 263040 1 0 $X=336110 $Y=258830
X1345 249 252 1 2 1089 XNR2D1BWP7T $T=184080 278720 0 0 $X=183790 $Y=278485
X1346 316 328 1 2 1135 XNR2D1BWP7T $T=236160 255200 0 0 $X=235870 $Y=254965
X1347 1134 363 1 2 1156 XNR2D1BWP7T $T=261360 278720 1 0 $X=261070 $Y=274510
X1348 1136 371 1 2 1153 XNR2D1BWP7T $T=264720 270880 1 0 $X=264430 $Y=266670
X1349 571 566 1 2 1257 XNR2D1BWP7T $T=404160 231680 0 0 $X=403870 $Y=231445
X1350 852 1 2 850 CKND0BWP7T $T=24480 255200 0 180 $X=22510 $Y=250990
X1351 854 1 2 952 CKND0BWP7T $T=84960 247360 0 0 $X=84670 $Y=247125
X1352 998 1 2 150 CKND0BWP7T $T=123600 247360 1 180 $X=121630 $Y=247125
X1353 202 1 2 206 CKND0BWP7T $T=155520 231680 0 0 $X=155230 $Y=231445
X1354 213 1 2 1056 CKND0BWP7T $T=171760 255200 0 180 $X=169790 $Y=250990
X1355 1128 1 2 318 CKND0BWP7T $T=263040 270880 1 0 $X=262750 $Y=266670
X1356 211 247 1 2 271 CKXOR2D0BWP7T $T=194160 294400 1 0 $X=193870 $Y=290190
X1357 1039 2 1040 1033 192 1034 1 AOI22D2BWP7T $T=157200 278720 1 180 $X=150190 $Y=278485
X1358 211 2 1040 1057 192 1045 1 AOI22D2BWP7T $T=163920 278720 1 0 $X=163630 $Y=274510
X1359 214 2 1045 1027 211 219 1 AOI22D2BWP7T $T=163920 286560 0 0 $X=163630 $Y=286325
X1360 1062 2 198 1069 197 1032 1 AOI22D2BWP7T $T=170640 278720 1 0 $X=170350 $Y=274510
X1361 1044 2 1045 1041 211 216 1 AOI22D2BWP7T $T=170640 286560 0 0 $X=170350 $Y=286325
X1362 1129 2 1115 329 324 320 1 AOI22D2BWP7T $T=233920 294400 1 0 $X=233630 $Y=290190
X1363 1159 2 1104 369 366 1132 1 AOI22D2BWP7T $T=261920 286560 1 0 $X=261630 $Y=282350
X1364 361 2 273 372 368 365 1 AOI22D2BWP7T $T=261920 294400 1 0 $X=261630 $Y=290190
X1365 337 2 284 385 366 380 1 AOI22D2BWP7T $T=268640 294400 1 0 $X=268350 $Y=290190
X1366 381 2 1157 399 1169 391 1 AOI22D2BWP7T $T=271440 278720 1 0 $X=271150 $Y=274510
X1367 381 2 334 405 1171 391 1 AOI22D2BWP7T $T=272560 263040 0 0 $X=272270 $Y=262805
X1368 381 2 393 390 1177 391 1 AOI22D2BWP7T $T=275360 270880 1 0 $X=275070 $Y=266670
X1369 381 2 319 438 429 391 1 AOI22D2BWP7T $T=298320 255200 0 0 $X=298030 $Y=254965
X1370 381 2 425 434 1192 391 1 AOI22D2BWP7T $T=298880 263040 1 0 $X=298590 $Y=258830
X1371 448 2 463 470 392 450 1 AOI22D2BWP7T $T=317360 286560 0 0 $X=317070 $Y=286325
X1372 1213 2 1104 482 366 486 1 AOI22D2BWP7T $T=335280 286560 1 0 $X=334990 $Y=282350
X1373 522 2 1230 1237 1233 527 1 AOI22D2BWP7T $T=373920 255200 1 0 $X=373630 $Y=250990
X1374 448 2 556 544 546 450 1 AOI22D2BWP7T $T=395200 294400 0 180 $X=388190 $Y=290190
X1375 448 2 595 590 583 450 1 AOI22D2BWP7T $T=428240 278720 0 180 $X=421230 $Y=274510
X1376 448 2 606 600 599 450 1 AOI22D2BWP7T $T=434400 270880 1 180 $X=427390 $Y=270645
X1377 448 2 618 621 484 450 1 AOI22D2BWP7T $T=441680 286560 0 180 $X=434670 $Y=282350
X1378 448 2 601 629 609 450 1 AOI22D2BWP7T $T=436080 278720 1 0 $X=435790 $Y=274510
X1379 448 2 310 631 1128 450 1 AOI22D2BWP7T $T=437760 270880 1 0 $X=437470 $Y=266670
X1380 1065 1062 1032 1064 1 2 MUX2ND0BWP7T $T=172880 278720 0 0 $X=172590 $Y=278485
X1381 1113 1128 318 1133 1 2 MUX2ND0BWP7T $T=233920 255200 1 0 $X=233630 $Y=250990
X1382 370 1169 1172 1167 1 2 MUX2ND0BWP7T $T=267520 255200 1 0 $X=267230 $Y=250990
X1383 397 1177 1181 402 1 2 MUX2ND0BWP7T $T=278160 239520 1 0 $X=277870 $Y=235310
X1384 464 439 1201 1202 1 2 MUX2ND0BWP7T $T=321840 247360 1 180 $X=317070 $Y=247125
X1385 1011 165 167 168 1014 2 1 AOI22D0BWP7T $T=132560 286560 1 0 $X=132270 $Y=282350
X1386 239 1070 1068 213 1056 2 1 AOI22D0BWP7T $T=182960 255200 0 180 $X=179310 $Y=250990
X1387 1089 1091 1080 1081 1061 2 1 AOI22D0BWP7T $T=189680 270880 0 0 $X=189390 $Y=270645
X1388 1156 1155 1134 340 349 2 1 AOI22D0BWP7T $T=259120 278720 1 180 $X=255470 $Y=278485
X1389 335 1204 458 381 391 2 1 AOI22D0BWP7T $T=320160 263040 0 180 $X=316510 $Y=258830
X1390 436 1205 456 448 450 2 1 AOI22D0BWP7T $T=320160 278720 0 180 $X=316510 $Y=274510
X1391 454 1203 462 381 391 2 1 AOI22D0BWP7T $T=317920 255200 1 0 $X=317630 $Y=250990
X1392 226 1066 258 2 1 1076 XNR3D0BWP7T $T=183520 263040 0 0 $X=183230 $Y=262805
X1393 1069 262 266 2 1 270 XNR3D0BWP7T $T=189680 278720 0 0 $X=189390 $Y=278485
X1394 887 1 2 149 CKBD0BWP7T $T=112400 286560 1 0 $X=112110 $Y=282350
X1395 187 1 2 1030 CKBD0BWP7T $T=148240 239520 1 0 $X=147950 $Y=235310
X1396 1046 1 2 1047 CKBD0BWP7T $T=163920 255200 0 0 $X=163630 $Y=254965
X1397 856 2 896 20 1 NR2D1BWP7T $T=60320 255200 0 180 $X=57790 $Y=250990
X1398 84 2 900 78 1 NR2D1BWP7T $T=71520 286560 1 180 $X=68990 $Y=286325
X1399 914 2 943 941 1 NR2D1BWP7T $T=82160 278720 1 180 $X=79630 $Y=278485
X1400 953 2 949 97 1 NR2D1BWP7T $T=84400 294400 1 0 $X=84110 $Y=290190
X1401 95 2 119 104 1 NR2D1BWP7T $T=95040 239520 1 0 $X=94750 $Y=235310
X1402 856 2 984 29 1 NR2D1BWP7T $T=107360 255200 0 180 $X=104830 $Y=250990
X1403 994 2 993 37 1 NR2D1BWP7T $T=114640 247360 0 180 $X=112110 $Y=243150
X1404 1002 2 1010 176 1 NR2D1BWP7T $T=142640 247360 1 180 $X=140110 $Y=247125
X1405 915 2 1007 5 1 NR2D1BWP7T $T=141520 263040 1 0 $X=141230 $Y=258830
X1406 435 2 1190 431 1 NR2D1BWP7T $T=306720 239520 0 180 $X=304190 $Y=235310
X1407 1207 2 1211 478 1 NR2D1BWP7T $T=333040 247360 0 0 $X=332750 $Y=247125
X1408 566 2 1258 431 1 NR2D1BWP7T $T=406400 239520 1 0 $X=406110 $Y=235310
X1409 1019 1020 163 178 1 2 AOI21D0BWP7T $T=144320 294400 0 180 $X=141230 $Y=290190
X1410 1141 1146 338 1145 1 2 AOI21D0BWP7T $T=251840 247360 1 0 $X=251550 $Y=243150
X1411 1140 1142 344 323 1 2 AOI21D0BWP7T $T=257440 255200 0 0 $X=257150 $Y=254965
X1412 1158 1160 1162 1165 1 2 AOI21D0BWP7T $T=260800 247360 1 0 $X=260510 $Y=243150
X1413 375 1170 351 323 1 2 AOI21D0BWP7T $T=270320 247360 1 180 $X=267230 $Y=247125
X1414 1175 1182 409 413 1 2 AOI21D0BWP7T $T=289920 278720 0 0 $X=289630 $Y=278485
X1415 430 1193 433 1197 1 2 AOI21D0BWP7T $T=303360 247360 1 0 $X=303070 $Y=243150
X1416 521 1238 532 323 1 2 AOI21D0BWP7T $T=379520 239520 0 0 $X=379230 $Y=239285
X1417 1255 1260 580 1259 1 2 AOI21D0BWP7T $T=419280 255200 1 180 $X=416190 $Y=254965
X1418 1256 1262 582 413 1 2 AOI21D0BWP7T $T=420960 239520 0 180 $X=417870 $Y=235310
X1419 865 22 9 12 2 1 863 NR4D1BWP7T $T=31200 270880 0 180 $X=25310 $Y=266670
X1420 875 876 9 26 2 1 863 NR4D1BWP7T $T=45760 270880 1 180 $X=39870 $Y=270645
X1421 925 73 920 904 2 1 69 NR4D1BWP7T $T=66480 286560 1 180 $X=60590 $Y=286325
X1422 72 910 78 885 2 1 882 NR4D1BWP7T $T=65360 255200 1 0 $X=65070 $Y=250990
X1423 956 93 94 100 2 1 104 NR4D1BWP7T $T=83840 231680 0 0 $X=83550 $Y=231445
X1424 964 96 91 80 2 1 882 NR4D1BWP7T $T=96720 247360 1 180 $X=90830 $Y=247125
X1425 959 110 7 960 2 1 966 NR4D1BWP7T $T=91680 270880 0 0 $X=91390 $Y=270645
X1426 970 84 879 906 2 1 891 NR4D1BWP7T $T=99520 255200 1 180 $X=93630 $Y=254965
X1427 133 125 974 962 2 1 914 NR4D1BWP7T $T=103440 278720 1 180 $X=97550 $Y=278485
X1428 140 84 127 989 2 1 991 NR4D1BWP7T $T=106240 255200 0 0 $X=105950 $Y=254965
X1429 995 148 146 143 2 1 139 NR4D1BWP7T $T=115200 231680 1 180 $X=109310 $Y=231445
X1430 1028 145 62 975 2 1 1016 NR4D1BWP7T $T=148800 263040 1 180 $X=142910 $Y=262805
X1431 68 2 928 54 881 20 1 AOI31D2BWP7T $T=61440 239520 0 0 $X=61150 $Y=239285
X1432 37 54 897 954 1 2 998 OA31D0BWP7T $T=127520 255200 0 180 $X=122750 $Y=250990
X1433 852 1 3 847 2 ND2D1BWP7T $T=24480 270880 0 0 $X=24190 $Y=270645
X1434 852 1 17 24 2 ND2D1BWP7T $T=26720 294400 1 0 $X=26430 $Y=290190
X1435 25 1 849 852 2 ND2D1BWP7T $T=29520 286560 0 180 $X=26990 $Y=282350
X1436 18 1 858 25 2 ND2D1BWP7T $T=31200 278720 1 180 $X=28670 $Y=278485
X1437 18 1 27 861 2 ND2D1BWP7T $T=28960 286560 0 0 $X=28670 $Y=286325
X1438 864 1 859 868 2 ND2D1BWP7T $T=37920 255200 1 0 $X=37630 $Y=250990
X1439 859 1 884 874 2 ND2D1BWP7T $T=42400 263040 1 0 $X=42110 $Y=258830
X1440 852 1 860 868 2 ND2D1BWP7T $T=45200 247360 1 0 $X=44910 $Y=243150
X1441 864 1 39 24 2 ND2D1BWP7T $T=45200 286560 0 0 $X=44910 $Y=286325
X1442 847 1 44 19 2 ND2D1BWP7T $T=52480 270880 1 180 $X=49950 $Y=270645
X1443 19 1 51 24 2 ND2D1BWP7T $T=53600 286560 0 180 $X=51070 $Y=282350
X1444 54 1 878 893 2 ND2D1BWP7T $T=54160 239520 1 180 $X=51630 $Y=239285
X1445 902 1 898 51 2 ND2D1BWP7T $T=55280 255200 1 180 $X=52750 $Y=254965
X1446 44 1 895 903 2 ND2D1BWP7T $T=53040 278720 1 0 $X=52750 $Y=274510
X1447 881 1 52 19 2 ND2D1BWP7T $T=56400 278720 1 180 $X=53870 $Y=278485
X1448 10 1 56 900 2 ND2D1BWP7T $T=58080 294400 0 180 $X=55550 $Y=290190
X1449 907 1 903 861 2 ND2D1BWP7T $T=58640 278720 1 180 $X=56110 $Y=278485
X1450 862 1 906 59 2 ND2D1BWP7T $T=56960 278720 1 0 $X=56670 $Y=274510
X1451 24 1 57 908 2 ND2D1BWP7T $T=56960 286560 1 0 $X=56670 $Y=282350
X1452 18 1 43 881 2 ND2D1BWP7T $T=58640 278720 0 0 $X=58350 $Y=278485
X1453 847 1 912 55 2 ND2D1BWP7T $T=59200 263040 0 0 $X=58910 $Y=262805
X1454 25 1 65 908 2 ND2D1BWP7T $T=61440 286560 0 180 $X=58910 $Y=282350
X1455 847 1 899 864 2 ND2D1BWP7T $T=59760 270880 0 0 $X=59470 $Y=270645
X1456 916 1 67 864 2 ND2D1BWP7T $T=63680 263040 1 180 $X=61150 $Y=262805
X1457 852 1 917 916 2 ND2D1BWP7T $T=62000 263040 1 0 $X=61710 $Y=258830
X1458 917 1 66 899 2 ND2D1BWP7T $T=64240 278720 0 180 $X=61710 $Y=274510
X1459 868 1 855 921 2 ND2D1BWP7T $T=62560 255200 0 0 $X=62270 $Y=254965
X1460 847 1 902 921 2 ND2D1BWP7T $T=64240 263040 1 0 $X=63950 $Y=258830
X1461 27 1 924 855 2 ND2D1BWP7T $T=67040 278720 1 180 $X=64510 $Y=278485
X1462 881 1 926 864 2 ND2D1BWP7T $T=67600 270880 1 180 $X=65070 $Y=270645
X1463 83 1 80 27 2 ND2D1BWP7T $T=69280 286560 0 180 $X=66750 $Y=282350
X1464 872 1 919 881 2 ND2D1BWP7T $T=70400 270880 0 180 $X=67870 $Y=266670
X1465 847 1 922 907 2 ND2D1BWP7T $T=73200 278720 0 180 $X=70670 $Y=274510
X1466 847 1 913 908 2 ND2D1BWP7T $T=83280 278720 0 180 $X=80750 $Y=274510
X1467 872 1 934 847 2 ND2D1BWP7T $T=86640 270880 0 180 $X=84110 $Y=266670
X1468 25 1 954 907 2 ND2D1BWP7T $T=85520 255200 0 0 $X=85230 $Y=254965
X1469 47 1 98 951 2 ND2D1BWP7T $T=85520 278720 1 0 $X=85230 $Y=274510
X1470 907 1 112 868 2 ND2D1BWP7T $T=87760 255200 0 0 $X=87470 $Y=254965
X1471 916 1 947 921 2 ND2D1BWP7T $T=91120 263040 0 180 $X=88590 $Y=258830
X1472 916 1 31 908 2 ND2D1BWP7T $T=91120 263040 1 180 $X=88590 $Y=262805
X1473 18 1 890 916 2 ND2D1BWP7T $T=91120 278720 0 180 $X=88590 $Y=274510
X1474 39 1 960 899 2 ND2D1BWP7T $T=93360 278720 0 180 $X=90830 $Y=274510
X1475 25 1 83 921 2 ND2D1BWP7T $T=91680 263040 1 0 $X=91390 $Y=258830
X1476 116 1 122 938 2 ND2D1BWP7T $T=95040 231680 0 0 $X=94750 $Y=231445
X1477 881 1 106 921 2 ND2D1BWP7T $T=97840 263040 1 180 $X=95310 $Y=262805
X1478 120 1 968 112 2 ND2D1BWP7T $T=98400 286560 1 180 $X=95870 $Y=286325
X1479 908 1 969 868 2 ND2D1BWP7T $T=101760 255200 0 180 $X=99230 $Y=250990
X1480 39 1 974 979 2 ND2D1BWP7T $T=100640 278720 1 0 $X=100350 $Y=274510
X1481 131 1 978 43 2 ND2D1BWP7T $T=104560 294400 0 180 $X=102030 $Y=290190
X1482 967 1 135 903 2 ND2D1BWP7T $T=107920 278720 1 180 $X=105390 $Y=278485
X1483 872 1 120 916 2 ND2D1BWP7T $T=124160 270880 1 180 $X=121630 $Y=270645
X1484 83 1 999 913 2 ND2D1BWP7T $T=121920 278720 1 0 $X=121630 $Y=274510
X1485 983 1 159 908 2 ND2D1BWP7T $T=131440 255200 0 180 $X=128910 $Y=250990
X1486 881 1 985 908 2 ND2D1BWP7T $T=134800 263040 1 180 $X=132270 $Y=262805
X1487 983 1 851 155 2 ND2D1BWP7T $T=137040 255200 1 180 $X=134510 $Y=254965
X1488 176 1 946 155 2 ND2D1BWP7T $T=140400 247360 1 180 $X=137870 $Y=247125
X1489 1002 1 973 176 2 ND2D1BWP7T $T=143760 255200 0 0 $X=143470 $Y=254965
X1490 849 1 3 848 2 853 856 OAI211D1BWP7T $T=22240 286560 1 0 $X=21950 $Y=282350
X1491 860 1 919 70 2 920 14 OAI211D1BWP7T $T=65360 247360 1 180 $X=61710 $Y=247125
X1492 860 1 919 70 2 937 14 OAI211D1BWP7T $T=69840 247360 0 0 $X=69550 $Y=247125
X1493 947 1 909 4 2 958 946 OAI211D1BWP7T $T=84960 263040 0 0 $X=84670 $Y=262805
X1494 111 1 59 973 2 124 29 OAI211D1BWP7T $T=98960 294400 1 0 $X=98670 $Y=290190
X1495 964 1 870 13 2 126 982 OAI211D1BWP7T $T=100640 247360 0 0 $X=100350 $Y=247125
X1496 874 1 992 973 2 166 915 OAI211D1BWP7T $T=136480 294400 0 180 $X=132830 $Y=290190
X1497 917 1 159 851 2 1016 14 OAI211D1BWP7T $T=137040 263040 0 180 $X=133390 $Y=258830
X1498 874 1 992 973 2 172 915 OAI211D1BWP7T $T=137600 294400 1 0 $X=137310 $Y=290190
X1499 1163 1 1151 354 2 357 336 OAI211D1BWP7T $T=261360 231680 1 180 $X=257710 $Y=231445
X1500 1155 1 355 323 2 1110 359 OAI211D1BWP7T $T=258560 294400 1 0 $X=258270 $Y=290190
X1501 1254 1 1253 1252 2 1245 336 OAI211D1BWP7T $T=405280 239520 1 180 $X=401630 $Y=239285
X1502 891 2 882 879 867 1 33 NR4D2BWP7T $T=51360 247360 1 180 $X=38190 $Y=247125
X1503 871 2 12 888 891 1 53 NR4D2BWP7T $T=40160 255200 1 0 $X=39870 $Y=250990
X1504 884 2 889 22 876 1 870 NR4D2BWP7T $T=45200 263040 0 0 $X=44910 $Y=262805
X1505 888 2 85 885 78 1 108 NR4D2BWP7T $T=92800 255200 0 180 $X=79630 $Y=250990
X1506 862 1 859 858 855 11 2 ND4D1BWP7T $T=27840 278720 0 180 $X=23630 $Y=274510
X1507 890 1 48 42 849 46 2 ND4D1BWP7T $T=51920 294400 0 180 $X=47710 $Y=290190
X1508 909 1 903 51 57 58 2 ND4D1BWP7T $T=60320 286560 1 180 $X=56110 $Y=286325
X1509 922 1 855 43 909 918 2 ND4D1BWP7T $T=64800 278720 1 180 $X=60590 $Y=278485
X1510 10 1 59 927 886 75 2 ND4D1BWP7T $T=64800 294400 1 0 $X=64510 $Y=290190
X1511 912 1 934 919 909 940 2 ND4D1BWP7T $T=69280 263040 0 0 $X=68990 $Y=262805
X1512 144 1 913 147 929 996 2 ND4D1BWP7T $T=111280 278720 0 0 $X=110990 $Y=278485
X1513 1002 1001 991 848 929 1 2 OAI31D1BWP7T $T=125840 255200 1 180 $X=121630 $Y=254965
X1514 940 125 1000 151 168 1 2 OAI31D1BWP7T $T=122480 286560 0 0 $X=122190 $Y=286325
X1515 924 932 158 965 163 1 2 OAI31D1BWP7T $T=127520 286560 1 0 $X=127230 $Y=282350
X1516 30 1 10 870 2 871 ND3D0BWP7T $T=42960 270880 0 180 $X=39870 $Y=266670
X1517 59 1 913 57 2 63 ND3D0BWP7T $T=62000 294400 0 180 $X=58910 $Y=290190
X1518 922 1 83 873 2 941 ND3D0BWP7T $T=70400 278720 0 0 $X=70110 $Y=278485
X1519 939 1 943 865 2 942 ND3D0BWP7T $T=82720 270880 0 180 $X=79630 $Y=266670
X1520 955 1 105 902 2 92 ND3D0BWP7T $T=87200 278720 1 180 $X=84110 $Y=278485
X1521 969 1 926 909 2 981 ND3D0BWP7T $T=100080 263040 0 0 $X=99790 $Y=262805
X1522 1002 1 907 155 2 955 ND3D0BWP7T $T=129200 255200 1 180 $X=126110 $Y=254965
X1523 896 1 2 889 879 911 910 NR4D0BWP7T $T=57520 255200 0 0 $X=57230 $Y=254965
X1524 936 1 2 879 99 101 103 NR4D0BWP7T $T=84960 286560 0 0 $X=84670 $Y=286325
X1525 932 1 2 972 971 121 99 NR4D0BWP7T $T=101760 286560 1 180 $X=98110 $Y=286325
X1526 846 4 2 6 1 NR2D2BWP7T $T=21120 239520 1 0 $X=20830 $Y=235310
X1527 850 5 2 15 1 NR2D2BWP7T $T=22800 255200 0 0 $X=22510 $Y=254965
X1528 897 915 2 933 1 NR2D2BWP7T $T=110720 239520 1 180 $X=106510 $Y=239285
X1529 855 3 877 880 2 1 40 AN4D1BWP7T $T=41840 278720 1 0 $X=41550 $Y=274510
X1530 886 43 874 849 2 1 880 AN4D1BWP7T $T=51360 286560 0 180 $X=47150 $Y=282350
X1531 875 1 2 883 BUFFD0BWP7T $T=42960 270880 1 0 $X=42670 $Y=266670
X1532 925 1 2 930 BUFFD0BWP7T $T=66480 286560 0 0 $X=66190 $Y=286325
X1533 893 868 901 37 898 2 1 AOI31D1BWP7T $T=53040 247360 0 0 $X=52750 $Y=247125
X1534 123 938 977 36 129 2 1 AOI31D1BWP7T $T=101200 239520 1 0 $X=100910 $Y=235310
X1535 31 1 859 849 28 869 2 ND4D0BWP7T $T=41840 286560 0 180 $X=38190 $Y=282350
X1536 862 1 39 47 51 45 2 ND4D0BWP7T $T=48560 286560 0 0 $X=48270 $Y=286325
X1537 44 1 865 40 900 904 2 ND4D0BWP7T $T=52480 286560 0 0 $X=52190 $Y=286325
X1538 31 1 83 927 928 87 2 ND4D0BWP7T $T=68720 294400 1 0 $X=68430 $Y=290190
X1539 65 1 922 34 947 953 2 ND4D0BWP7T $T=81040 286560 1 0 $X=80750 $Y=282350
X1540 105 1 934 899 922 113 2 ND4D0BWP7T $T=89440 278720 0 0 $X=89150 $Y=278485
X1541 31 1 10 947 961 962 2 ND4D0BWP7T $T=92240 263040 0 0 $X=91950 $Y=262805
X1542 31 1 115 943 117 965 2 ND4D0BWP7T $T=93360 286560 1 0 $X=93070 $Y=282350
X1543 131 1 976 926 43 972 2 ND4D0BWP7T $T=104000 286560 0 180 $X=100350 $Y=282350
X1544 954 1 988 959 886 141 2 ND4D0BWP7T $T=111280 278720 1 180 $X=107630 $Y=278485
X1545 985 1 106 34 108 989 2 ND4D0BWP7T $T=114080 263040 1 180 $X=110430 $Y=262805
X1546 955 1 934 1004 987 1011 2 ND4D0BWP7T $T=124160 278720 0 0 $X=123870 $Y=278485
X1547 990 1 957 149 1012 1013 2 ND4D0BWP7T $T=132000 278720 1 0 $X=131710 $Y=274510
X1548 967 1 1015 1006 1012 1014 2 ND4D0BWP7T $T=134800 270880 0 0 $X=134510 $Y=270645
X1549 970 1 175 108 1012 1019 2 ND4D0BWP7T $T=138720 278720 1 0 $X=138430 $Y=274510
X1550 887 2 86 98 153 1004 1 INR4D0BWP7T $T=129200 294400 0 180 $X=124430 $Y=290190
X1551 917 2 1007 958 174 1015 1 INR4D0BWP7T $T=142640 270880 0 180 $X=137870 $Y=266670
X1552 876 1 9 869 887 2 NR3D1BWP7T $T=41840 286560 1 0 $X=41550 $Y=282350
X1553 22 1 80 918 81 2 NR3D1BWP7T $T=70960 278720 0 180 $X=66190 $Y=274510
X1554 130 1 894 985 136 890 2 IND4D0BWP7T $T=104000 278720 1 0 $X=103710 $Y=274510
X1555 46 1 53 928 944 949 2 IND4D1BWP7T $T=79920 294400 1 0 $X=79630 $Y=290190
X1556 884 1 959 42 975 47 2 IND4D1BWP7T $T=89440 270880 1 0 $X=89150 $Y=266670
X1557 142 1 883 42 137 976 2 IND4D1BWP7T $T=110720 263040 1 180 $X=105950 $Y=262805
X1558 905 2 50 41 32 1 36 NR4D3BWP7T $T=57520 231680 1 180 $X=41550 $Y=231445
X1559 853 35 7 873 866 1 2 INR4D1BWP7T $T=44640 286560 1 180 $X=37630 $Y=286325
X1560 15 867 895 49 899 1 2 INR4D1BWP7T $T=48000 270880 1 0 $X=47710 $Y=266670
X1561 135 971 968 987 131 1 2 INR4D1BWP7T $T=110720 286560 1 180 $X=103710 $Y=286325
X1562 130 110 974 990 83 1 2 INR4D1BWP7T $T=114080 270880 1 180 $X=107070 $Y=270645
X1563 102 134 978 992 913 1 2 INR4D1BWP7T $T=108480 294400 1 0 $X=108190 $Y=290190
X1564 76 923 1 82 938 2 INR3D1BWP7T $T=66480 231680 0 0 $X=66190 $Y=231445
X1565 848 2 8 1 851 NR2XD1BWP7T $T=23360 263040 1 0 $X=23070 $Y=258830
X1566 13 2 21 1 846 NR2XD1BWP7T $T=26160 239520 1 0 $X=25870 $Y=235310
X1567 857 2 867 1 4 NR2XD1BWP7T $T=38480 239520 0 0 $X=38190 $Y=239285
X1568 20 2 61 1 54 NR2XD1BWP7T $T=56960 239520 0 0 $X=56670 $Y=239285
X1569 70 2 910 1 931 NR2XD1BWP7T $T=65920 247360 0 0 $X=65630 $Y=247125
X1570 897 2 78 1 4 NR2XD1BWP7T $T=83840 239520 1 180 $X=79630 $Y=239285
X1571 70 2 91 1 4 NR2XD1BWP7T $T=81040 247360 1 0 $X=80750 $Y=243150
X1572 931 2 96 1 5 NR2XD1BWP7T $T=84400 239520 0 0 $X=84110 $Y=239285
X1573 37 2 921 1 854 NR2XD1BWP7T $T=93360 247360 0 180 $X=89150 $Y=243150
X1574 13 2 145 1 946 NR2XD1BWP7T $T=110160 247360 0 0 $X=109870 $Y=247125
X1575 176 2 983 1 171 NR2XD1BWP7T $T=143200 255200 1 180 $X=138990 $Y=254965
X1576 516 2 514 1 431 NR2XD1BWP7T $T=365520 239520 0 180 $X=361310 $Y=235310
X1577 71 1 923 74 2 IND2D1BWP7T $T=63680 231680 0 0 $X=63390 $Y=231445
X1578 876 1 77 67 2 IND2D1BWP7T $T=69280 263040 1 180 $X=66190 $Y=262805
X1579 22 1 932 919 2 IND2D1BWP7T $T=67600 270880 0 0 $X=67310 $Y=270645
X1580 127 1 966 929 2 IND2D1BWP7T $T=105680 270880 0 180 $X=102590 $Y=266670
X1581 77 8 885 933 2 1 935 OR4XD1BWP7T $T=68160 255200 0 0 $X=67870 $Y=254965
X1582 104 128 132 114 2 1 986 OR4XD1BWP7T $T=102880 231680 0 0 $X=102590 $Y=231445
X1583 874 2 889 898 64 62 1 INR4D2BWP7T $T=46880 263040 1 0 $X=46590 $Y=258830
X1584 874 1 992 973 2 915 160 OAI211D0BWP7T $T=133120 294400 0 180 $X=129470 $Y=290190
X1585 1000 1 1020 1022 2 186 1025 OAI211D0BWP7T $T=144880 286560 0 0 $X=144590 $Y=286325
X1586 315 1 1131 323 2 1133 1121 OAI211D0BWP7T $T=236160 239520 0 0 $X=235870 $Y=239285
X1587 849 1 3 856 23 848 2 OAI211D2BWP7T $T=22240 286560 0 0 $X=21950 $Y=286325
X1588 859 1 855 5 26 854 2 OAI211D2BWP7T $T=24480 255200 1 0 $X=24190 $Y=250990
X1589 1018 1 1017 181 184 182 2 OAI211D2BWP7T $T=141520 239520 1 0 $X=141230 $Y=235310
X1590 1018 1 1017 181 188 182 2 OAI211D2BWP7T $T=143760 239520 0 0 $X=143470 $Y=239285
X1591 1021 1 1029 186 199 1028 2 OAI211D2BWP7T $T=148240 286560 0 0 $X=147950 $Y=286325
X1592 187 1 190 194 200 191 2 OAI211D2BWP7T $T=148800 231680 0 0 $X=148510 $Y=231445
X1593 1030 1 190 194 196 191 2 OAI211D2BWP7T $T=151040 239520 1 0 $X=150750 $Y=235310
X1594 1148 1 1147 336 333 1137 2 OAI211D2BWP7T $T=256320 255200 0 180 $X=249870 $Y=250990
X1595 18 1 24 866 2 CKND2D0BWP7T $T=28960 294400 1 0 $X=28670 $Y=290190
X1596 872 868 1007 997 1 2 142 AO211D0BWP7T $T=130320 263040 1 180 $X=126110 $Y=262805
X1597 1010 872 137 999 1 2 1005 AO211D0BWP7T $T=130320 270880 1 180 $X=126110 $Y=270645
X1598 312 480 465 476 1 2 1209 AO211D0BWP7T $T=336960 231680 1 180 $X=332750 $Y=231445
X1599 936 2 937 957 952 916 1 AOI211D2BWP7T $T=81040 263040 1 0 $X=80750 $Y=258830
X1600 850 2 9 857 1 NR2D3BWP7T $T=21120 247360 0 0 $X=20830 $Y=247125
X1601 854 2 852 20 1 NR2D3BWP7T $T=23360 247360 1 0 $X=23070 $Y=243150
X1602 14 2 19 20 1 NR2D3BWP7T $T=25600 231680 0 0 $X=25310 $Y=231445
X1603 878 2 864 20 1 NR2D3BWP7T $T=45760 239520 0 180 $X=40430 $Y=235310
X1604 897 2 85 931 1 NR2D3BWP7T $T=68160 239520 0 0 $X=67870 $Y=239285
X1605 13 2 84 5 1 NR2D3BWP7T $T=97840 239520 0 0 $X=97550 $Y=239285
X1606 52 863 890 1 2 ND2D2BWP7T $T=50240 278720 0 0 $X=49950 $Y=278485
X1607 61 29 893 1 2 ND2D2BWP7T $T=61440 247360 0 180 $X=57230 $Y=243150
X1608 1001 897 983 1 2 ND2D2BWP7T $T=125280 247360 0 0 $X=124990 $Y=247125
X1609 868 42 18 1 2 ND2D2BWP7T $T=129760 263040 1 0 $X=129470 $Y=258830
X1610 941 1 2 89 879 948 NR3D0BWP7T $T=80480 286560 0 0 $X=80190 $Y=286325
X1611 924 1 2 984 933 961 NR3D0BWP7T $T=107360 263040 0 180 $X=104270 $Y=258830
X1612 110 1 2 885 997 1006 NR3D0BWP7T $T=124160 263040 1 0 $X=123870 $Y=258830
X1613 497 1216 1 1217 492 2 AOI21D1BWP7T $T=346480 239520 0 180 $X=342830 $Y=235310
X1614 591 1261 1 1264 592 2 AOI21D1BWP7T $T=424880 286560 1 180 $X=421230 $Y=286325
X1615 30 969 127 934 2 1 ND3D2BWP7T $T=97280 270880 0 0 $X=96990 $Y=270645
X1616 171 176 963 1001 2 1 ND3D2BWP7T $T=142640 247360 0 180 $X=137310 $Y=243150
X1617 39 899 926 10 69 1 2 ND4D2BWP7T $T=93360 286560 0 180 $X=85790 $Y=282350
X1618 163 1 161 945 96 981 2 OAI31D2BWP7T $T=132000 278720 0 180 $X=124990 $Y=274510
X1619 167 1 1021 996 980 118 2 OAI31D2BWP7T $T=146000 278720 1 180 $X=138990 $Y=278485
X1620 111 1 106 42 2 35 ND3D1BWP7T $T=92800 294400 0 180 $X=89150 $Y=290190
X1621 31 1 874 948 2 118 ND3D1BWP7T $T=92800 286560 0 0 $X=92510 $Y=286325
X1622 969 1 144 120 2 130 ND3D1BWP7T $T=111280 278720 1 0 $X=110990 $Y=274510
X1623 102 2 867 952 1 951 847 AOI211D1BWP7T $T=87200 270880 1 180 $X=83550 $Y=270645
X1624 906 2 879 907 1 979 983 AOI211D1BWP7T $T=102320 255200 0 0 $X=102030 $Y=254965
X1625 1160 2 341 351 1 1151 312 AOI211D1BWP7T $T=259120 239520 1 180 $X=255470 $Y=239285
X1626 1194 2 1190 428 1 1189 312 AOI211D1BWP7T $T=304480 278720 0 180 $X=300830 $Y=274510
X1627 1211 2 323 1207 1 1208 478 AOI211D1BWP7T $T=336960 247360 0 0 $X=336670 $Y=247125
X1628 536 2 514 521 1 520 312 AOI211D1BWP7T $T=377280 231680 1 180 $X=373630 $Y=231445
X1629 1260 2 1258 1255 1 1253 312 AOI211D1BWP7T $T=419280 239520 1 180 $X=415630 $Y=239285
X1630 584 2 1258 1257 1 579 312 AOI211D1BWP7T $T=420400 231680 1 180 $X=416750 $Y=231445
X1631 926 2 927 15 1 INR2D1BWP7T $T=72080 286560 0 180 $X=68990 $Y=282350
X1650 613 460 2 1 CKBD2BWP7T $T=434960 239520 1 180 $X=431310 $Y=239285
X1651 1 2 ICV_21 $T=26720 270880 0 0 $X=26430 $Y=270645
X1652 1 2 ICV_21 $T=93360 247360 1 0 $X=93070 $Y=243150
X1653 1 2 ICV_21 $T=135360 286560 0 0 $X=135070 $Y=286325
X1654 1 2 ICV_21 $T=194720 286560 1 0 $X=194430 $Y=282350
X1655 1 2 ICV_21 $T=227200 270880 0 0 $X=226910 $Y=270645
X1656 1 2 ICV_21 $T=278720 239520 0 0 $X=278430 $Y=239285
X1657 1 2 ICV_21 $T=278720 270880 0 0 $X=278430 $Y=270645
X1658 1 2 ICV_21 $T=298880 270880 0 0 $X=298590 $Y=270645
X1659 1 2 ICV_21 $T=310080 247360 0 0 $X=309790 $Y=247125
X1660 1 2 ICV_21 $T=320720 231680 0 0 $X=320430 $Y=231445
X1661 1 2 ICV_21 $T=338080 278720 1 0 $X=337790 $Y=274510
X1662 1 2 ICV_21 $T=362720 239520 0 0 $X=362430 $Y=239285
X1663 1 2 ICV_21 $T=362720 263040 0 0 $X=362430 $Y=262805
X1664 1 2 ICV_21 $T=380640 255200 1 0 $X=380350 $Y=250990
X1665 1 2 ICV_21 $T=396880 231680 0 0 $X=396590 $Y=231445
X1666 1 2 ICV_21 $T=413120 263040 1 0 $X=412830 $Y=258830
X1667 1 2 ICV_21 $T=419280 255200 0 0 $X=418990 $Y=254965
X1668 1 2 ICV_21 $T=422080 278720 0 0 $X=421790 $Y=278485
X1669 1 2 ICV_21 $T=429360 255200 0 0 $X=429070 $Y=254965
X1670 1 2 ICV_21 $T=429920 294400 1 0 $X=429630 $Y=290190
X1671 1 2 ICV_21 $T=446720 294400 1 0 $X=446430 $Y=290190
X1676 268 1118 287 1282 2 1 306 DFCND1BWP7T $T=220480 286560 0 0 $X=220190 $Y=286325
X1677 268 1119 257 1283 2 1 300 DFCND1BWP7T $T=222720 255200 0 0 $X=222430 $Y=254965
X1678 268 322 257 1284 2 1 307 DFCND1BWP7T $T=240640 231680 1 180 $X=227470 $Y=231445
X1679 268 346 257 360 2 1 1143 DFCND1BWP7T $T=251840 263040 0 0 $X=251550 $Y=262805
X1680 468 1215 282 1285 2 1 1199 DFCND1BWP7T $T=352080 255200 0 180 $X=338910 $Y=250990
X1681 468 1219 282 1286 2 1 339 DFCND1BWP7T $T=352080 270880 0 180 $X=338910 $Y=266670
X1682 468 1218 282 505 2 1 507 DFCND1BWP7T $T=346480 278720 0 0 $X=346190 $Y=278485
X1683 468 1248 282 1287 2 1 542 DFCND1BWP7T $T=400800 255200 1 180 $X=387630 $Y=254965
X1684 468 1242 282 1288 2 1 554 DFCND1BWP7T $T=388480 278720 0 0 $X=388190 $Y=278485
X1685 997 1 2 984 993 988 916 AOI211XD0BWP7T $T=115200 255200 1 180 $X=111550 $Y=254965
X1686 162 1 2 977 157 1009 156 AOI211XD0BWP7T $T=131440 239520 0 180 $X=127790 $Y=235310
X1687 1146 1 2 341 1140 1147 312 AOI211XD0BWP7T $T=255200 247360 1 180 $X=251550 $Y=247125
X1688 356 1 2 341 1135 1152 312 AOI211XD0BWP7T $T=260800 247360 1 180 $X=257150 $Y=247125
X1689 1208 1 2 465 1207 459 312 AOI211XD0BWP7T $T=323520 239520 1 180 $X=319870 $Y=239285
X1690 268 1120 257 313 1130 1 2 DFCND2BWP7T $T=223280 247360 0 0 $X=222990 $Y=247125
X1691 268 1122 287 320 1129 1 2 DFCND2BWP7T $T=225520 286560 1 0 $X=225230 $Y=282350
X1692 268 1144 257 1159 1132 1 2 DFCND2BWP7T $T=249040 263040 1 0 $X=248750 $Y=258830
X1693 468 494 282 481 479 1 2 DFCND2BWP7T $T=348720 294400 0 180 $X=333870 $Y=290190
X1694 468 1220 282 486 1213 1 2 DFCND2BWP7T $T=352080 286560 1 180 $X=337230 $Y=286325
X1695 468 1224 282 496 493 1 2 DFCND2BWP7T $T=359920 270880 1 180 $X=345070 $Y=270645
X1696 468 1221 282 510 512 1 2 DFCND2BWP7T $T=347600 255200 0 0 $X=347310 $Y=254965
X1697 468 1229 282 1223 1222 1 2 DFCND2BWP7T $T=366080 247360 1 180 $X=351230 $Y=247125
X1698 468 1240 282 555 553 1 2 DFCND2BWP7T $T=382320 231680 0 0 $X=382030 $Y=231445
X1699 468 1244 552 569 1251 1 2 DFCND2BWP7T $T=390720 278720 1 0 $X=390430 $Y=274510
X1700 919 1 68 897 13 2 OAI21D2BWP7T $T=70960 239520 0 180 $X=65630 $Y=235310
X1701 967 1 888 848 856 2 OAI21D2BWP7T $T=97840 255200 0 180 $X=92510 $Y=250990
X1702 926 1 102 29 963 2 OAI21D2BWP7T $T=98400 263040 1 0 $X=98110 $Y=258830
X1703 1152 1 358 323 1166 2 OAI21D2BWP7T $T=265840 247360 1 180 $X=260510 $Y=247125
X1704 421 1 1107 418 1185 2 OAI21D2BWP7T $T=298320 239520 0 180 $X=292990 $Y=235310
X1705 424 1 1108 376 1188 2 OAI21D2BWP7T $T=299440 247360 1 180 $X=294110 $Y=247125
X1706 1210 1 483 323 1212 2 OAI21D2BWP7T $T=331920 255200 0 0 $X=331630 $Y=254965
X1707 535 1 1123 418 1232 2 OAI21D2BWP7T $T=381760 270880 1 180 $X=376430 $Y=270645
X1708 539 1 529 515 537 2 OAI21D2BWP7T $T=385120 294400 0 180 $X=379790 $Y=290190
X1709 1179 395 1 1116 386 2 IOA21D1BWP7T $T=279840 286560 0 180 $X=276190 $Y=282350
X1710 1200 427 1 423 1189 2 IOA21D1BWP7T $T=302800 278720 1 180 $X=299150 $Y=278485
X1711 1263 549 1 1112 585 2 IOA21D1BWP7T $T=423760 263040 0 180 $X=420110 $Y=258830
X1712 524 528 1234 1236 531 1 2 533 AO221D1BWP7T $T=375600 278720 1 0 $X=375310 $Y=274510
X1713 508 649 1276 1278 531 1 2 662 AO221D1BWP7T $T=461840 239520 0 0 $X=461550 $Y=239285
X1714 317 656 1280 1281 531 1 2 663 AO221D1BWP7T $T=461840 278720 1 0 $X=461550 $Y=274510
X1715 268 291 257 1289 2 1 1085 DFCND0BWP7T $T=220480 247360 0 180 $X=207310 $Y=243150
X1716 268 1125 257 1290 2 1 1117 DFCND0BWP7T $T=235600 263040 0 180 $X=222430 $Y=258830
X1717 268 1126 287 1291 2 1 1114 DFCND0BWP7T $T=236160 278720 0 180 $X=222990 $Y=274510
X1718 268 325 257 1292 2 1 308 DFCND0BWP7T $T=241200 239520 0 180 $X=228030 $Y=235310
X1719 268 1149 257 1139 2 1 330 DFCND0BWP7T $T=261360 239520 0 180 $X=248190 $Y=235310
X1720 468 1206 282 1293 2 1 1198 DFCND0BWP7T $T=324080 263040 1 180 $X=310910 $Y=262805
X1721 468 1241 282 1230 2 1 1233 DFCND0BWP7T $T=390720 247360 0 180 $X=377550 $Y=243150
X1722 468 1243 552 1249 2 1 1250 DFCND0BWP7T $T=388480 286560 1 0 $X=388190 $Y=282350
X1723 383 376 373 379 364 1139 2 1150 1 OA222D0BWP7T $T=274240 239520 0 180 $X=267790 $Y=235310
X1724 1231 418 501 1230 387 496 2 1228 1 OA222D0BWP7T $T=366080 270880 0 180 $X=359630 $Y=266670
X1725 1234 515 501 499 387 505 2 1227 1 OA222D0BWP7T $T=384000 286560 1 180 $X=377550 $Y=286325
X1726 543 515 501 568 387 1249 2 1246 1 OA222D0BWP7T $T=405280 286560 1 180 $X=398830 $Y=286325
X1727 574 515 501 570 387 567 2 1247 1 OA222D0BWP7T $T=406400 294400 0 180 $X=399950 $Y=290190
X1728 578 515 501 567 387 588 2 1265 1 OA222D0BWP7T $T=416480 294400 1 0 $X=416190 $Y=290190
X1729 11 2 38 1 894 892 896 AOI211XD1BWP7T $T=46320 278720 1 0 $X=46030 $Y=274510
X1730 1193 2 1190 1 437 312 430 AOI211XD1BWP7T $T=308960 239520 1 180 $X=301950 $Y=239285
X1731 229 233 1 2 INVD6BWP7T $T=172880 231680 0 0 $X=172590 $Y=231445
X1732 376 384 1 373 1159 364 367 2 1161 OAI222D2BWP7T $T=274240 231680 1 180 $X=263870 $Y=231445
X1733 418 498 1 501 1223 387 509 2 1226 OAI222D2BWP7T $T=349840 247360 1 0 $X=349550 $Y=243150
X1734 515 519 1 501 481 387 506 2 504 OAI222D2BWP7T $T=364960 294400 0 180 $X=354590 $Y=290190
X1735 515 517 1 501 486 387 1223 2 1220 OAI222D2BWP7T $T=366080 286560 1 180 $X=355710 $Y=286325
X1736 418 518 1 501 510 387 481 2 1221 OAI222D2BWP7T $T=366640 263040 0 180 $X=356270 $Y=258830
X1737 491 1 2 431 INVD5BWP7T $T=345360 231680 0 0 $X=345070 $Y=231445
X1738 13 2 1 963 876 NR2D2P5BWP7T $T=91680 239520 0 0 $X=91390 $Y=239285
X1739 973 2 1 155 24 NR2D2P5BWP7T $T=144320 278720 1 0 $X=144030 $Y=274510
X1740 986 122 152 1003 154 1 2 OAI31D0BWP7T $T=123600 231680 0 0 $X=123310 $Y=231445
X1741 864 25 22 2 1 CKAN2D2BWP7T $T=31200 263040 0 180 $X=26990 $Y=258830
X1742 109 2 95 923 88 1 NR3D2BWP7T $T=90560 239520 0 180 $X=80190 $Y=235310
X1743 171 946 856 1 2 OR2D2BWP7T $T=137600 247360 1 180 $X=133390 $Y=247125
X1744 274 275 279 1 2 OR2D2BWP7T $T=206480 239520 1 0 $X=206190 $Y=235310
X1745 852 10 16 1 2 ND2D1P5BWP7T $T=23920 263040 0 0 $X=23630 $Y=262805
X1746 864 874 16 1 2 ND2D1P5BWP7T $T=43520 263040 1 180 $X=39310 $Y=262805
X1747 20 915 55 1 2 ND2D1P5BWP7T $T=64240 239520 0 180 $X=60030 $Y=235310
X1748 892 854 54 1 2 ND2D1P5BWP7T $T=123600 239520 0 0 $X=123310 $Y=239285
X1749 994 14 892 1 2 ND2D1P5BWP7T $T=128640 239520 0 0 $X=128350 $Y=239285
X1750 1010 846 1001 1 2 ND2D1P5BWP7T $T=135920 239520 0 0 $X=135630 $Y=239285
X1751 27 886 876 1 2 INR2XD1BWP7T $T=48560 278720 1 180 $X=43790 $Y=278485
X1752 18 848 1 2 INVD1P5BWP7T $T=23920 278720 1 180 $X=21390 $Y=278485
X1753 336 349 1 2 CKND6BWP7T $T=295520 278720 1 0 $X=295230 $Y=274510
X1754 623 1 1162 654 647 1279 2 1277 OAI221D2BWP7T $T=469680 255200 1 180 $X=460430 $Y=254965
X1755 1 2 ICV_23 $T=35120 247360 1 0 $X=34830 $Y=243150
X1756 1 2 ICV_23 $T=35120 255200 0 0 $X=34830 $Y=254965
X1757 1 2 ICV_23 $T=245120 247360 0 0 $X=244830 $Y=247125
X1758 1 2 ICV_23 $T=245120 263040 0 0 $X=244830 $Y=262805
X1759 1 2 ICV_23 $T=306720 239520 1 0 $X=306430 $Y=235310
X1760 1 2 ICV_23 $T=310640 286560 1 0 $X=310350 $Y=282350
X1761 1 2 ICV_23 $T=329120 286560 0 0 $X=328830 $Y=286325
X1762 1 2 ICV_23 $T=384000 286560 0 0 $X=383710 $Y=286325
X1763 1 2 ICV_23 $T=390720 247360 1 0 $X=390430 $Y=243150
X1764 1 2 ICV_23 $T=395760 270880 0 0 $X=395470 $Y=270645
X1765 1 2 ICV_23 $T=405280 239520 0 0 $X=404990 $Y=239285
X1766 1 2 ICV_23 $T=405280 278720 1 0 $X=404990 $Y=274510
X1767 1 2 ICV_23 $T=405280 286560 0 0 $X=404990 $Y=286325
X1768 1 2 ICV_23 $T=413120 278720 1 0 $X=412830 $Y=274510
X1769 1 2 ICV_23 $T=413120 286560 0 0 $X=412830 $Y=286325
X1770 1 2 ICV_23 $T=429920 239520 1 0 $X=429630 $Y=235310
X1771 1 2 ICV_23 $T=447280 255200 1 0 $X=446990 $Y=250990
X1772 1 2 ICV_23 $T=447280 263040 0 0 $X=446990 $Y=262805
X1773 1 2 ICV_23 $T=455120 239520 0 0 $X=454830 $Y=239285
X1774 1 2 ICV_23 $T=455120 278720 1 0 $X=454830 $Y=274510
X1775 212 217 223 225 1 2 1059 AO22D0BWP7T $T=166720 270880 0 0 $X=166430 $Y=270645
X1776 412 2 391 1 CKND10BWP7T $T=292160 231680 0 0 $X=291870 $Y=231445
X1777 171 155 176 2 5 1 ND3D3BWP7T $T=146000 255200 0 0 $X=145710 $Y=254965
X1778 171 155 1031 881 1 2 AN3D2BWP7T $T=152160 270880 1 180 $X=147390 $Y=270645
X1779 895 1 901 912 914 2 IND3D2BWP7T $T=56400 270880 1 0 $X=56110 $Y=266670
X1780 864 1 861 34 2 CKND2D2BWP7T $T=41840 294400 1 0 $X=41550 $Y=290190
X1798 236 534 1231 1239 531 540 1 2 AO221D2BWP7T $T=378960 263040 0 0 $X=378670 $Y=262805
X1799 643 582 1275 1274 531 658 1 2 AO221D2BWP7T $T=459040 239520 1 0 $X=458750 $Y=235310
X1800 1 2 ICV_26 $T=236160 278720 1 0 $X=235870 $Y=274510
X1801 1 2 ICV_26 $T=264720 263040 0 0 $X=264430 $Y=262805
X1802 1 2 ICV_26 $T=287120 286560 0 0 $X=286830 $Y=286325
X1803 1 2 ICV_26 $T=294400 239520 0 0 $X=294110 $Y=239285
X1804 1 2 ICV_26 $T=320160 263040 1 0 $X=319870 $Y=258830
X1805 1 2 ICV_26 $T=320160 286560 1 0 $X=319870 $Y=282350
X1806 1 2 ICV_26 $T=336960 231680 0 0 $X=336670 $Y=231445
X1807 1 2 ICV_26 $T=352080 270880 1 0 $X=351790 $Y=266670
X1808 1 2 ICV_26 $T=362160 255200 0 0 $X=361870 $Y=254965
X1809 1 2 ICV_26 $T=381760 270880 0 0 $X=381470 $Y=270645
X1810 1 2 ICV_26 $T=389600 270880 1 0 $X=389310 $Y=266670
X1811 1 2 ICV_26 $T=392960 255200 1 0 $X=392670 $Y=250990
X1812 1 2 ICV_26 $T=398560 239520 1 0 $X=398270 $Y=235310
X1813 1 2 ICV_26 $T=419840 270880 0 0 $X=419550 $Y=270645
X1814 1 2 ICV_26 $T=428240 278720 1 0 $X=427950 $Y=274510
X1815 1 2 ICV_26 $T=431600 247360 1 0 $X=431310 $Y=243150
X1816 1 2 ICV_26 $T=455120 270880 0 0 $X=454830 $Y=270645
X1817 1 2 ICV_27 $T=20000 239520 0 0 $X=19710 $Y=239285
X1818 1 2 ICV_27 $T=20000 270880 0 0 $X=19710 $Y=270645
X1819 1 2 ICV_27 $T=34000 247360 0 0 $X=33710 $Y=247125
X1820 1 2 ICV_27 $T=76000 255200 0 0 $X=75710 $Y=254965
X1821 1 2 ICV_27 $T=160000 247360 1 0 $X=159710 $Y=243150
X1822 1 2 ICV_27 $T=160000 270880 0 0 $X=159710 $Y=270645
X1823 1 2 ICV_27 $T=202000 231680 0 0 $X=201710 $Y=231445
X1824 1 2 ICV_27 $T=202000 239520 1 0 $X=201710 $Y=235310
X1825 1 2 ICV_27 $T=244000 231680 0 0 $X=243710 $Y=231445
X1826 1 2 ICV_27 $T=244000 239520 1 0 $X=243710 $Y=235310
X1827 1 2 ICV_27 $T=244000 239520 0 0 $X=243710 $Y=239285
X1828 1 2 ICV_27 $T=244000 270880 0 0 $X=243710 $Y=270645
X1829 1 2 ICV_27 $T=244000 278720 0 0 $X=243710 $Y=278485
X1830 1 2 ICV_27 $T=286000 294400 1 0 $X=285710 $Y=290190
X1831 1 2 ICV_27 $T=328000 239520 1 0 $X=327710 $Y=235310
X1832 1 2 ICV_27 $T=370000 270880 1 0 $X=369710 $Y=266670
X1833 1 2 ICV_27 $T=412000 247360 0 0 $X=411710 $Y=247125
X1834 1 2 ICV_27 $T=412000 255200 0 0 $X=411710 $Y=254965
X1835 1 2 ICV_27 $T=412000 294400 1 0 $X=411710 $Y=290190
X1836 1 2 ICV_27 $T=454000 255200 1 0 $X=453710 $Y=250990
X1837 1237 1 336 525 1235 413 2 OAI22D2BWP7T $T=382880 255200 1 180 $X=375870 $Y=254965
X1838 336 1196 1194 413 1195 2 1 OAI22D0BWP7T $T=307840 278720 0 180 $X=304190 $Y=274510
X1839 209 218 1 2 BUFFD4BWP7T $T=163920 231680 0 0 $X=163630 $Y=231445
X1840 54 2 892 37 1 18 NR3D3BWP7T $T=154400 255200 0 180 $X=142350 $Y=250990
X1841 164 1008 177 169 1 179 2 ND4D4BWP7T $T=133120 231680 0 0 $X=132830 $Y=231445
X1842 868 61 980 29 2 982 1 IOA22D2BWP7T $T=100640 247360 1 0 $X=100350 $Y=243150
X1843 897 16 1 2 CKND8BWP7T $T=53600 239520 0 180 $X=46590 $Y=235310
X1844 19 25 885 1 2 AN2D2BWP7T $T=43520 255200 0 0 $X=43230 $Y=254965
X1845 21 860 7 1 2 IND2D2BWP7T $T=28960 239520 1 180 $X=24190 $Y=239285
.ENDS
***************************************
.SUBCKT NR2XD3BWP7T A2 VDD A1 VSS ZN
** N=6 EP=5 IP=0 FDC=20
M0 VSS A2 ZN VSS N L=1.8e-07 W=6e-07 $X=820 $Y=345 $D=0
M1 ZN A2 VSS VSS N L=1.8e-07 W=6e-07 $X=1540 $Y=345 $D=0
M2 VSS A2 ZN VSS N L=1.8e-07 W=6e-07 $X=2260 $Y=345 $D=0
M3 ZN A2 VSS VSS N L=1.8e-07 W=6e-07 $X=2980 $Y=345 $D=0
M4 VSS A2 ZN VSS N L=1.8e-07 W=6e-07 $X=3700 $Y=345 $D=0
M5 ZN A1 VSS VSS N L=1.8e-07 W=6e-07 $X=4420 $Y=345 $D=0
M6 VSS A1 ZN VSS N L=1.8e-07 W=6e-07 $X=5140 $Y=345 $D=0
M7 ZN A1 VSS VSS N L=1.8e-07 W=6e-07 $X=5860 $Y=345 $D=0
M8 VSS A1 ZN VSS N L=1.8e-07 W=6e-07 $X=6580 $Y=345 $D=0
M9 ZN A1 VSS VSS N L=1.8e-07 W=6e-07 $X=7300 $Y=345 $D=0
M10 6 A2 VDD VDD P L=1.8e-07 W=1.14e-06 $X=820 $Y=2435 $D=16
M11 VDD A2 6 VDD P L=1.8e-07 W=1.77e-06 $X=1540 $Y=1805 $D=16
M12 6 A2 VDD VDD P L=1.8e-07 W=1.77e-06 $X=2260 $Y=1805 $D=16
M13 VDD A2 6 VDD P L=1.8e-07 W=1.77e-06 $X=2980 $Y=1805 $D=16
M14 6 A2 VDD VDD P L=1.8e-07 W=1.77e-06 $X=3700 $Y=1805 $D=16
M15 ZN A1 6 VDD P L=1.8e-07 W=1.77e-06 $X=4420 $Y=1805 $D=16
M16 6 A1 ZN VDD P L=1.8e-07 W=1.77e-06 $X=5140 $Y=1805 $D=16
M17 ZN A1 6 VDD P L=1.8e-07 W=1.77e-06 $X=5860 $Y=1805 $D=16
M18 6 A1 ZN VDD P L=1.8e-07 W=1.77e-06 $X=6580 $Y=1805 $D=16
M19 ZN A1 6 VDD P L=1.8e-07 W=1.14e-06 $X=7300 $Y=2435 $D=16
.ENDS
***************************************
.SUBCKT EDFCND2BWP7T E D CP CDN QN Q VSS VDD
** N=25 EP=8 IP=0 FDC=42
M0 VSS E 9 VSS N L=1.8e-07 W=5e-07 $X=620 $Y=505 $D=0
M1 19 D VSS VSS N L=1.8e-07 W=5.7e-07 $X=1380 $Y=775 $D=0
M2 12 E 19 VSS N L=1.8e-07 W=5.7e-07 $X=1810 $Y=775 $D=0
M3 20 9 12 VSS N L=1.8e-07 W=4.2e-07 $X=2570 $Y=650 $D=0
M4 VSS 16 20 VSS N L=1.8e-07 W=4.2e-07 $X=3000 $Y=650 $D=0
M5 VSS CP 10 VSS N L=1.8e-07 W=5e-07 $X=4260 $Y=980 $D=0
M6 11 10 VSS VSS N L=1.8e-07 W=5e-07 $X=4865 $Y=980 $D=0
M7 14 10 12 VSS N L=1.8e-07 W=7.4e-07 $X=6285 $Y=575 $D=0
M8 21 11 14 VSS N L=1.8e-07 W=4.2e-07 $X=7115 $Y=895 $D=0
M9 22 CDN 21 VSS N L=1.8e-07 W=4.2e-07 $X=7575 $Y=895 $D=0
M10 VSS 15 22 VSS N L=1.8e-07 W=4.2e-07 $X=8035 $Y=895 $D=0
M11 15 14 VSS VSS N L=1.8e-07 W=5.4e-07 $X=8895 $Y=775 $D=0
M12 17 11 15 VSS N L=1.8e-07 W=9.1e-07 $X=9770 $Y=405 $D=0
M13 16 10 17 VSS N L=1.8e-07 W=4.2e-07 $X=10535 $Y=895 $D=0
M14 VSS 18 16 VSS N L=1.8e-07 W=1e-06 $X=12170 $Y=345 $D=0
M15 23 CDN VSS VSS N L=1.8e-07 W=9.3e-07 $X=12950 $Y=345 $D=0
M16 18 17 23 VSS N L=1.8e-07 W=1e-06 $X=13640 $Y=345 $D=0
M17 QN 16 VSS VSS N L=1.8e-07 W=1e-06 $X=15520 $Y=345 $D=0
M18 VSS 16 QN VSS N L=1.8e-07 W=1e-06 $X=16240 $Y=345 $D=0
M19 Q 18 VSS VSS N L=1.8e-07 W=1e-06 $X=16960 $Y=345 $D=0
M20 VSS 18 Q VSS N L=1.8e-07 W=1e-06 $X=17680 $Y=345 $D=0
M21 VDD E 9 VDD P L=1.8e-07 W=6.85e-07 $X=620 $Y=2830 $D=16
M22 24 D VDD VDD P L=1.8e-07 W=7.5e-07 $X=1380 $Y=2395 $D=16
M23 12 9 24 VDD P L=1.8e-07 W=7.5e-07 $X=1810 $Y=2395 $D=16
M24 25 E 12 VDD P L=1.8e-07 W=4.2e-07 $X=2530 $Y=2725 $D=16
M25 VDD 16 25 VDD P L=1.8e-07 W=4.2e-07 $X=2960 $Y=2725 $D=16
M26 VDD CP 10 VDD P L=1.8e-07 W=6.85e-07 $X=4260 $Y=2345 $D=16
M27 11 10 VDD VDD P L=1.8e-07 W=6.85e-07 $X=4870 $Y=2345 $D=16
M28 14 11 12 VDD P L=1.8e-07 W=7.8e-07 $X=6290 $Y=2345 $D=16
M29 13 10 14 VDD P L=1.8e-07 W=4.2e-07 $X=7145 $Y=2345 $D=16
M30 VDD CDN 13 VDD P L=1.8e-07 W=4.2e-07 $X=7865 $Y=2345 $D=16
M31 13 15 VDD VDD P L=1.8e-07 W=4.2e-07 $X=8465 $Y=2345 $D=16
M32 15 14 VDD VDD P L=1.8e-07 W=6.2e-07 $X=9735 $Y=2175 $D=16
M33 17 10 15 VDD P L=1.8e-07 W=6.2e-07 $X=10535 $Y=2175 $D=16
M34 16 11 17 VDD P L=1.8e-07 W=4.2e-07 $X=11450 $Y=2205 $D=16
M35 VDD 18 16 VDD P L=1.8e-07 W=1.37e-06 $X=12170 $Y=2205 $D=16
M36 18 CDN VDD VDD P L=1.8e-07 W=4.2e-07 $X=12950 $Y=2350 $D=16
M37 VDD 17 18 VDD P L=1.8e-07 W=1.37e-06 $X=14800 $Y=2205 $D=16
M38 QN 16 VDD VDD P L=1.8e-07 W=1.37e-06 $X=15520 $Y=2205 $D=16
M39 VDD 16 QN VDD P L=1.8e-07 W=1.37e-06 $X=16240 $Y=2205 $D=16
M40 Q 18 VDD VDD P L=1.8e-07 W=1.37e-06 $X=16960 $Y=2205 $D=16
M41 VDD 18 Q VDD P L=1.8e-07 W=1.37e-06 $X=17680 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT NR4D4BWP7T A4 VDD A3 A2 A1 ZN VSS
** N=10 EP=7 IP=0 FDC=56
M0 ZN A4 VSS VSS N L=1.8e-07 W=5.7e-07 $X=820 $Y=345 $D=0
M1 VSS A4 ZN VSS N L=1.8e-07 W=5.7e-07 $X=1545 $Y=345 $D=0
M2 ZN A4 VSS VSS N L=1.8e-07 W=5.7e-07 $X=2265 $Y=345 $D=0
M3 VSS A4 ZN VSS N L=1.8e-07 W=5.7e-07 $X=2985 $Y=345 $D=0
M4 ZN A4 VSS VSS N L=1.8e-07 W=5.7e-07 $X=3705 $Y=345 $D=0
M5 VSS A4 ZN VSS N L=1.8e-07 W=5.7e-07 $X=4425 $Y=345 $D=0
M6 ZN A4 VSS VSS N L=1.8e-07 W=5.7e-07 $X=5145 $Y=345 $D=0
M7 VSS A3 ZN VSS N L=1.8e-07 W=5.7e-07 $X=5865 $Y=345 $D=0
M8 ZN A3 VSS VSS N L=1.8e-07 W=5.7e-07 $X=6585 $Y=345 $D=0
M9 VSS A3 ZN VSS N L=1.8e-07 W=5.7e-07 $X=7305 $Y=345 $D=0
M10 ZN A3 VSS VSS N L=1.8e-07 W=5.7e-07 $X=8025 $Y=345 $D=0
M11 VSS A3 ZN VSS N L=1.8e-07 W=5.7e-07 $X=8745 $Y=345 $D=0
M12 ZN A3 VSS VSS N L=1.8e-07 W=5.7e-07 $X=9465 $Y=345 $D=0
M13 VSS A3 ZN VSS N L=1.8e-07 W=5.7e-07 $X=10185 $Y=345 $D=0
M14 ZN A2 VSS VSS N L=1.8e-07 W=5.7e-07 $X=10905 $Y=345 $D=0
M15 VSS A2 ZN VSS N L=1.8e-07 W=5.7e-07 $X=11625 $Y=345 $D=0
M16 ZN A2 VSS VSS N L=1.8e-07 W=5.7e-07 $X=12345 $Y=345 $D=0
M17 VSS A2 ZN VSS N L=1.8e-07 W=5.7e-07 $X=13065 $Y=345 $D=0
M18 ZN A2 VSS VSS N L=1.8e-07 W=5.7e-07 $X=13785 $Y=345 $D=0
M19 VSS A2 ZN VSS N L=1.8e-07 W=5.7e-07 $X=14505 $Y=345 $D=0
M20 ZN A2 VSS VSS N L=1.8e-07 W=5.7e-07 $X=15225 $Y=345 $D=0
M21 VSS A1 ZN VSS N L=1.8e-07 W=5.7e-07 $X=15945 $Y=345 $D=0
M22 ZN A1 VSS VSS N L=1.8e-07 W=5.7e-07 $X=16665 $Y=345 $D=0
M23 VSS A1 ZN VSS N L=1.8e-07 W=5.7e-07 $X=17385 $Y=345 $D=0
M24 ZN A1 VSS VSS N L=1.8e-07 W=5.7e-07 $X=18105 $Y=345 $D=0
M25 VSS A1 ZN VSS N L=1.8e-07 W=5.7e-07 $X=18825 $Y=345 $D=0
M26 ZN A1 VSS VSS N L=1.8e-07 W=5.7e-07 $X=19545 $Y=345 $D=0
M27 VSS A1 ZN VSS N L=1.8e-07 W=5.7e-07 $X=20265 $Y=345 $D=0
M28 8 A4 VDD VDD P L=1.8e-07 W=1.36e-06 $X=820 $Y=2215 $D=16
M29 VDD A4 8 VDD P L=1.8e-07 W=1.6e-06 $X=1545 $Y=1975 $D=16
M30 8 A4 VDD VDD P L=1.8e-07 W=1.6e-06 $X=2265 $Y=1975 $D=16
M31 VDD A4 8 VDD P L=1.8e-07 W=1.6e-06 $X=2985 $Y=1975 $D=16
M32 8 A4 VDD VDD P L=1.8e-07 W=1.6e-06 $X=3705 $Y=1975 $D=16
M33 VDD A4 8 VDD P L=1.8e-07 W=1.6e-06 $X=4425 $Y=1975 $D=16
M34 8 A4 VDD VDD P L=1.8e-07 W=1.6e-06 $X=5145 $Y=1975 $D=16
M35 9 A3 8 VDD P L=1.8e-07 W=1.6e-06 $X=5865 $Y=1975 $D=16
M36 8 A3 9 VDD P L=1.8e-07 W=1.6e-06 $X=6585 $Y=1975 $D=16
M37 9 A3 8 VDD P L=1.8e-07 W=1.6e-06 $X=7305 $Y=1975 $D=16
M38 8 A3 9 VDD P L=1.8e-07 W=1.6e-06 $X=8025 $Y=1975 $D=16
M39 9 A3 8 VDD P L=1.8e-07 W=1.6e-06 $X=8745 $Y=1975 $D=16
M40 8 A3 9 VDD P L=1.8e-07 W=1.6e-06 $X=9465 $Y=1975 $D=16
M41 9 A3 8 VDD P L=1.8e-07 W=1.6e-06 $X=10185 $Y=1975 $D=16
M42 10 A2 9 VDD P L=1.8e-07 W=1.6e-06 $X=10905 $Y=1975 $D=16
M43 9 A2 10 VDD P L=1.8e-07 W=1.6e-06 $X=11625 $Y=1975 $D=16
M44 10 A2 9 VDD P L=1.8e-07 W=1.6e-06 $X=12345 $Y=1975 $D=16
M45 9 A2 10 VDD P L=1.8e-07 W=1.6e-06 $X=13065 $Y=1975 $D=16
M46 10 A2 9 VDD P L=1.8e-07 W=1.6e-06 $X=13785 $Y=1975 $D=16
M47 9 A2 10 VDD P L=1.8e-07 W=1.6e-06 $X=14505 $Y=1975 $D=16
M48 10 A2 9 VDD P L=1.8e-07 W=1.6e-06 $X=15225 $Y=1975 $D=16
M49 ZN A1 10 VDD P L=1.8e-07 W=1.6e-06 $X=15945 $Y=1975 $D=16
M50 10 A1 ZN VDD P L=1.8e-07 W=1.6e-06 $X=16665 $Y=1975 $D=16
M51 ZN A1 10 VDD P L=1.8e-07 W=1.6e-06 $X=17385 $Y=1975 $D=16
M52 10 A1 ZN VDD P L=1.8e-07 W=1.6e-06 $X=18105 $Y=1975 $D=16
M53 ZN A1 10 VDD P L=1.8e-07 W=1.6e-06 $X=18825 $Y=1975 $D=16
M54 10 A1 ZN VDD P L=1.8e-07 W=1.6e-06 $X=19545 $Y=1975 $D=16
M55 ZN A1 10 VDD P L=1.8e-07 W=1.36e-06 $X=20265 $Y=2215 $D=16
.ENDS
***************************************
.SUBCKT OR2D0BWP7T A1 VSS A2 VDD Z
** N=7 EP=5 IP=0 FDC=6
M0 6 A1 VSS VSS N L=1.8e-07 W=5e-07 $X=660 $Y=800 $D=0
M1 VSS A2 6 VSS N L=1.8e-07 W=5e-07 $X=1380 $Y=800 $D=0
M2 Z 6 VSS VSS N L=1.8e-07 W=5e-07 $X=2000 $Y=800 $D=0
M3 7 A1 6 VDD P L=1.8e-07 W=6.85e-07 $X=660 $Y=2885 $D=16
M4 VDD A2 7 VDD P L=1.8e-07 W=6.85e-07 $X=1200 $Y=2885 $D=16
M5 Z 6 VDD VDD P L=1.8e-07 W=6.85e-07 $X=2000 $Y=2885 $D=16
.ENDS
***************************************
.SUBCKT IIND4D0BWP7T A1 VSS B1 B2 ZN VDD A2
** N=12 EP=7 IP=0 FDC=12
M0 VSS A1 8 VSS N L=1.8e-07 W=4.2e-07 $X=620 $Y=460 $D=0
M1 10 8 ZN VSS N L=1.8e-07 W=5e-07 $X=1940 $Y=840 $D=0
M2 11 B1 10 VSS N L=1.8e-07 W=5e-07 $X=2490 $Y=840 $D=0
M3 12 B2 11 VSS N L=1.8e-07 W=5e-07 $X=3040 $Y=840 $D=0
M4 VSS 9 12 VSS N L=1.8e-07 W=5e-07 $X=3590 $Y=840 $D=0
M5 9 A2 VSS VSS N L=1.8e-07 W=4.2e-07 $X=4240 $Y=605 $D=0
M6 VDD A1 8 VDD P L=1.8e-07 W=4.2e-07 $X=620 $Y=2825 $D=16
M7 ZN 8 VDD VDD P L=1.8e-07 W=6.85e-07 $X=1345 $Y=2825 $D=16
M8 VDD B1 ZN VDD P L=1.8e-07 W=6.85e-07 $X=2065 $Y=2825 $D=16
M9 ZN B2 VDD VDD P L=1.8e-07 W=6.85e-07 $X=2800 $Y=2825 $D=16
M10 VDD 9 ZN VDD P L=1.8e-07 W=6.85e-07 $X=3520 $Y=2825 $D=16
M11 9 A2 VDD VDD P L=1.8e-07 W=4.2e-07 $X=4240 $Y=2825 $D=16
.ENDS
***************************************
.SUBCKT IINR4D1BWP7T B2 B1 ZN A2 VDD A1 VSS
** N=15 EP=7 IP=0 FDC=16
M0 ZN B1 VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS B2 ZN VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 ZN 9 VSS VSS N L=1.8e-07 W=7e-07 $X=3230 $Y=345 $D=0
M3 VSS 10 ZN VSS N L=1.8e-07 W=1e-06 $X=3950 $Y=345 $D=0
M4 VSS A2 9 VSS N L=1.8e-07 W=5e-07 $X=5640 $Y=460 $D=0
M5 10 A1 VSS VSS N L=1.8e-07 W=5e-07 $X=6470 $Y=460 $D=0
M6 11 B1 8 VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M7 VDD B2 11 VDD P L=1.8e-07 W=1.37e-06 $X=1100 $Y=2205 $D=16
M8 12 B2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=1820 $Y=2205 $D=16
M9 13 B1 12 VDD P L=1.8e-07 W=1.37e-06 $X=2350 $Y=2205 $D=16
M10 14 9 13 VDD P L=1.8e-07 W=1.37e-06 $X=2880 $Y=2205 $D=16
M11 ZN 10 14 VDD P L=1.8e-07 W=1.37e-06 $X=3410 $Y=2205 $D=16
M12 15 10 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4130 $Y=2205 $D=16
M13 8 9 15 VDD P L=1.8e-07 W=1.37e-06 $X=4580 $Y=2205 $D=16
M14 VDD A2 9 VDD P L=1.8e-07 W=6.85e-07 $X=5880 $Y=2260 $D=16
M15 10 A1 VDD VDD P L=1.8e-07 W=6.85e-07 $X=6480 $Y=2260 $D=16
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480
+ 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 498 499 500 501
+ 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521
+ 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541
+ 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561
+ 562 563 564 565 566 567
** N=972 EP=566 IP=3602 FDC=4951
M0 970 834 1 1 N L=1.8e-07 W=5e-07 $X=129270 $Y=216460 $D=0
M1 971 144 970 1 N L=1.8e-07 W=5e-07 $X=129990 $Y=216460 $D=0
M2 851 843 971 1 N L=1.8e-07 W=5e-07 $X=130710 $Y=216460 $D=0
M3 972 130 851 1 N L=1.8e-07 W=5e-07 $X=131435 $Y=216460 $D=0
M4 1 144 972 1 N L=1.8e-07 W=5e-07 $X=132155 $Y=216460 $D=0
M5 853 851 1 1 N L=1.8e-07 W=5e-07 $X=133440 $Y=216460 $D=0
M6 850 834 851 2 P L=1.8e-07 W=6.85e-07 $X=129270 $Y=218550 $D=16
M7 851 144 850 2 P L=1.8e-07 W=6.85e-07 $X=129995 $Y=218550 $D=16
M8 850 843 851 2 P L=1.8e-07 W=6.85e-07 $X=130715 $Y=218550 $D=16
M9 2 130 850 2 P L=1.8e-07 W=6.85e-07 $X=131435 $Y=218550 $D=16
M10 850 144 2 2 P L=1.8e-07 W=6.85e-07 $X=132155 $Y=218340 $D=16
M11 853 851 2 2 P L=1.8e-07 W=6.85e-07 $X=133440 $Y=218805 $D=16
X90 1 506 ANTENNABWP7T $T=470800 223840 0 180 $X=469390 $Y=219630
X91 1 558 ANTENNABWP7T $T=470800 200320 0 0 $X=470510 $Y=200085
X92 1 543 ANTENNABWP7T $T=471920 208160 0 180 $X=470510 $Y=203950
X93 1 389 ANTENNABWP7T $T=470800 208160 0 0 $X=470510 $Y=207925
X94 1 396 ANTENNABWP7T $T=471920 216000 0 180 $X=470510 $Y=211790
X95 1 369 ANTENNABWP7T $T=470800 216000 0 0 $X=470510 $Y=215765
X96 1 520 ANTENNABWP7T $T=471920 223840 0 180 $X=470510 $Y=219630
X97 1 559 ANTENNABWP7T $T=470800 223840 0 0 $X=470510 $Y=223605
X98 1 560 ANTENNABWP7T $T=471920 231680 0 180 $X=470510 $Y=227470
X99 1 555 ANTENNABWP7T $T=471920 200320 0 0 $X=471630 $Y=200085
X100 1 564 ANTENNABWP7T $T=473040 208160 0 180 $X=471630 $Y=203950
X101 1 563 ANTENNABWP7T $T=471920 208160 0 0 $X=471630 $Y=207925
X102 1 498 ANTENNABWP7T $T=473040 216000 0 180 $X=471630 $Y=211790
X103 1 562 ANTENNABWP7T $T=471920 216000 0 0 $X=471630 $Y=215765
X104 1 539 ANTENNABWP7T $T=473040 223840 0 180 $X=471630 $Y=219630
X105 1 531 ANTENNABWP7T $T=471920 223840 0 0 $X=471630 $Y=223605
X106 1 509 ANTENNABWP7T $T=473040 231680 0 180 $X=471630 $Y=227470
X107 1 557 ANTENNABWP7T $T=473040 200320 0 0 $X=472750 $Y=200085
X108 1 565 ANTENNABWP7T $T=474160 208160 0 180 $X=472750 $Y=203950
X109 1 447 ANTENNABWP7T $T=473040 208160 0 0 $X=472750 $Y=207925
X110 1 458 ANTENNABWP7T $T=474160 216000 0 180 $X=472750 $Y=211790
X111 1 533 ANTENNABWP7T $T=473040 216000 0 0 $X=472750 $Y=215765
X112 1 566 ANTENNABWP7T $T=474160 223840 0 180 $X=472750 $Y=219630
X113 1 449 ANTENNABWP7T $T=473040 223840 0 0 $X=472750 $Y=223605
X114 1 567 ANTENNABWP7T $T=474160 231680 0 180 $X=472750 $Y=227470
X176 841 1 2 160 CKBD1BWP7T $T=137600 231680 1 0 $X=137310 $Y=227470
X177 257 1 2 891 CKBD1BWP7T $T=216560 208160 1 0 $X=216270 $Y=203950
X178 222 1 2 261 CKBD1BWP7T $T=219360 200320 0 0 $X=219070 $Y=200085
X179 337 1 2 889 CKBD1BWP7T $T=277600 208160 1 180 $X=275070 $Y=207925
X180 920 1 2 355 CKBD1BWP7T $T=294400 216000 1 180 $X=291870 $Y=215765
X181 369 1 2 366 CKBD1BWP7T $T=298880 223840 1 180 $X=296350 $Y=223605
X182 389 1 2 925 CKBD1BWP7T $T=323520 200320 1 180 $X=320990 $Y=200085
X183 533 1 2 532 CKBD1BWP7T $T=451200 208160 1 180 $X=448670 $Y=207925
X184 22 1 2 775 INVD0BWP7T $T=29520 231680 0 180 $X=27550 $Y=227470
X185 26 1 2 28 INVD0BWP7T $T=29520 216000 1 0 $X=29230 $Y=211790
X186 13 1 2 779 INVD0BWP7T $T=29520 216000 0 0 $X=29230 $Y=215765
X187 52 1 2 780 INVD0BWP7T $T=55280 208160 0 180 $X=53310 $Y=203950
X188 37 1 2 54 INVD0BWP7T $T=56960 208160 0 180 $X=54990 $Y=203950
X189 796 1 2 805 INVD0BWP7T $T=71520 223840 0 0 $X=71230 $Y=223605
X190 69 1 2 86 INVD0BWP7T $T=82160 231680 1 0 $X=81870 $Y=227470
X191 814 1 2 830 INVD0BWP7T $T=103440 216000 1 0 $X=103150 $Y=211790
X192 123 1 2 838 INVD0BWP7T $T=111280 200320 0 0 $X=110990 $Y=200085
X193 108 1 2 139 INVD0BWP7T $T=128640 231680 0 180 $X=126670 $Y=227470
X194 853 1 2 153 INVD0BWP7T $T=136480 231680 0 180 $X=134510 $Y=227470
X195 177 1 2 857 INVD0BWP7T $T=152720 231680 0 180 $X=150750 $Y=227470
X196 166 1 2 859 INVD0BWP7T $T=156640 231680 0 180 $X=154670 $Y=227470
X197 185 1 2 864 INVD0BWP7T $T=165040 208160 0 0 $X=164750 $Y=207925
X198 881 1 2 875 INVD0BWP7T $T=188000 216000 0 180 $X=186030 $Y=211790
X199 885 1 2 241 INVD0BWP7T $T=197520 208160 1 0 $X=197230 $Y=203950
X200 274 1 2 900 INVD0BWP7T $T=233360 231680 0 180 $X=231390 $Y=227470
X201 909 1 2 308 INVD0BWP7T $T=260800 223840 0 180 $X=258830 $Y=219630
X202 911 1 2 913 INVD0BWP7T $T=261360 208160 0 0 $X=261070 $Y=207925
X203 912 1 2 319 INVD0BWP7T $T=263600 200320 0 0 $X=263310 $Y=200085
X204 360 1 2 916 INVD0BWP7T $T=292720 216000 0 180 $X=290750 $Y=211790
X205 366 1 2 921 INVD0BWP7T $T=294960 223840 0 0 $X=294670 $Y=223605
X206 385 1 2 930 INVD0BWP7T $T=308960 223840 1 0 $X=308670 $Y=219630
X207 896 1 2 933 INVD0BWP7T $T=315680 231680 1 0 $X=315390 $Y=227470
X208 428 1 2 943 INVD0BWP7T $T=354320 223840 0 0 $X=354030 $Y=223605
X209 453 1 2 949 INVD0BWP7T $T=376720 216000 0 180 $X=374750 $Y=211790
X210 454 1 2 455 INVD0BWP7T $T=375600 200320 0 0 $X=375310 $Y=200085
X211 952 1 2 953 INVD0BWP7T $T=386240 223840 1 180 $X=384270 $Y=223605
X212 381 1 2 528 INVD0BWP7T $T=446160 231680 0 180 $X=444190 $Y=227470
X213 532 1 2 963 INVD0BWP7T $T=447840 208160 0 180 $X=445870 $Y=203950
X214 458 1 2 964 INVD0BWP7T $T=448960 216000 0 0 $X=448670 $Y=215765
X215 535 1 2 966 INVD0BWP7T $T=458480 216000 1 0 $X=458190 $Y=211790
X216 537 1 2 965 INVD0BWP7T $T=459600 223840 1 0 $X=459310 $Y=219630
X217 539 1 2 967 INVD0BWP7T $T=460720 231680 1 0 $X=460430 $Y=227470
X218 170 174 1 2 BUFFD1P5BWP7T $T=146560 200320 0 0 $X=146270 $Y=200085
X219 907 303 1 2 BUFFD1P5BWP7T $T=254640 208160 1 0 $X=254350 $Y=203950
X220 244 358 1 2 BUFFD1P5BWP7T $T=289920 223840 0 0 $X=289630 $Y=223605
X221 499 464 1 2 BUFFD1P5BWP7T $T=420400 216000 1 180 $X=417310 $Y=215765
X222 506 504 1 2 BUFFD1P5BWP7T $T=429920 216000 1 180 $X=426830 $Y=215765
X223 509 508 1 2 BUFFD1P5BWP7T $T=431600 216000 0 180 $X=428510 $Y=211790
X224 520 516 1 2 BUFFD1P5BWP7T $T=438880 208160 1 180 $X=435790 $Y=207925
X225 521 394 1 2 BUFFD1P5BWP7T $T=439440 216000 1 180 $X=436350 $Y=215765
X226 523 336 1 2 BUFFD1P5BWP7T $T=442800 208160 0 180 $X=439710 $Y=203950
X227 530 526 1 2 BUFFD1P5BWP7T $T=446160 208160 1 180 $X=443070 $Y=207925
X228 531 522 1 2 BUFFD1P5BWP7T $T=447280 216000 1 180 $X=444190 $Y=215765
X229 534 381 1 2 BUFFD1P5BWP7T $T=451200 223840 1 180 $X=448110 $Y=223605
X230 543 515 1 2 BUFFD1P5BWP7T $T=465200 216000 0 180 $X=462110 $Y=211790
X231 555 551 1 2 BUFFD1P5BWP7T $T=469680 223840 0 180 $X=466590 $Y=219630
X232 556 552 1 2 BUFFD1P5BWP7T $T=470800 216000 0 180 $X=467710 $Y=211790
X233 557 553 1 2 BUFFD1P5BWP7T $T=470800 231680 0 180 $X=467710 $Y=227470
X234 524 1 2 529 INVD3BWP7T $T=442240 216000 1 0 $X=441950 $Y=211790
X235 542 1 2 545 INVD3BWP7T $T=463520 208160 0 0 $X=463230 $Y=207925
X236 548 1 2 554 INVD3BWP7T $T=465760 200320 0 0 $X=465470 $Y=200085
X273 338 525 525 338 936 1 2 MAOI22D2BWP7T $T=445040 223840 0 180 $X=438590 $Y=219630
X274 787 1 2 44 BUFFD1BWP7T $T=49680 216000 0 0 $X=49390 $Y=215765
X275 826 1 2 834 BUFFD1BWP7T $T=106240 223840 1 0 $X=105950 $Y=219630
X276 836 1 2 856 BUFFD1BWP7T $T=142080 216000 0 0 $X=141790 $Y=215765
X277 847 1 2 167 BUFFD1BWP7T $T=144880 216000 0 0 $X=144590 $Y=215765
X278 872 1 2 870 BUFFD1BWP7T $T=176800 208160 1 0 $X=176510 $Y=203950
X279 887 1 2 242 BUFFD1BWP7T $T=196960 223840 0 0 $X=196670 $Y=223605
X280 371 1 2 370 BUFFD1BWP7T $T=299440 200320 1 180 $X=296910 $Y=200085
X281 922 1 2 373 BUFFD1BWP7T $T=302240 231680 0 180 $X=299710 $Y=227470
X282 923 1 2 380 BUFFD1BWP7T $T=302240 208160 1 0 $X=301950 $Y=203950
X283 926 1 2 388 BUFFD1BWP7T $T=305600 200320 0 0 $X=305310 $Y=200085
X284 892 1 2 406 BUFFD1BWP7T $T=319600 208160 0 0 $X=319310 $Y=207925
X285 410 1 2 408 BUFFD1BWP7T $T=324080 208160 0 180 $X=321550 $Y=203950
X286 452 1 2 451 BUFFD1BWP7T $T=376160 223840 1 180 $X=373630 $Y=223605
X287 962 1 2 519 BUFFD1BWP7T $T=434960 231680 1 0 $X=434670 $Y=227470
X288 1 2 DCAP4BWP7T $T=55280 200320 0 0 $X=54990 $Y=200085
X289 1 2 DCAP4BWP7T $T=94480 216000 0 0 $X=94190 $Y=215765
X290 1 2 DCAP4BWP7T $T=123600 208160 0 0 $X=123310 $Y=207925
X291 1 2 DCAP4BWP7T $T=138160 216000 1 0 $X=137870 $Y=211790
X292 1 2 DCAP4BWP7T $T=140400 223840 0 0 $X=140110 $Y=223605
X293 1 2 DCAP4BWP7T $T=157760 200320 0 0 $X=157470 $Y=200085
X294 1 2 DCAP4BWP7T $T=157760 223840 1 0 $X=157470 $Y=219630
X295 1 2 DCAP4BWP7T $T=241760 208160 1 0 $X=241470 $Y=203950
X296 1 2 DCAP4BWP7T $T=263600 216000 1 0 $X=263310 $Y=211790
X297 1 2 DCAP4BWP7T $T=319600 208160 1 0 $X=319310 $Y=203950
X298 1 2 DCAP4BWP7T $T=357680 200320 0 0 $X=357390 $Y=200085
X299 1 2 DCAP4BWP7T $T=392960 223840 1 0 $X=392670 $Y=219630
X300 1 2 DCAP4BWP7T $T=398560 216000 0 0 $X=398270 $Y=215765
X301 1 2 ICV_3 $T=21120 216000 0 0 $X=20830 $Y=215765
X302 1 2 ICV_3 $T=21120 223840 1 0 $X=20830 $Y=219630
X303 1 2 ICV_3 $T=31200 216000 1 0 $X=30910 $Y=211790
X304 1 2 ICV_3 $T=51920 216000 0 0 $X=51630 $Y=215765
X305 1 2 ICV_3 $T=92800 200320 0 0 $X=92510 $Y=200085
X306 1 2 ICV_3 $T=93920 208160 1 0 $X=93630 $Y=203950
X307 1 2 ICV_3 $T=115200 200320 0 0 $X=114910 $Y=200085
X308 1 2 ICV_3 $T=115200 216000 1 0 $X=114910 $Y=211790
X309 1 2 ICV_3 $T=115200 216000 0 0 $X=114910 $Y=215765
X310 1 2 ICV_3 $T=119120 200320 0 0 $X=118830 $Y=200085
X311 1 2 ICV_3 $T=119120 208160 1 0 $X=118830 $Y=203950
X312 1 2 ICV_3 $T=119120 223840 0 0 $X=118830 $Y=223605
X313 1 2 ICV_3 $T=125840 216000 0 0 $X=125550 $Y=215765
X314 1 2 ICV_3 $T=129760 208160 1 0 $X=129470 $Y=203950
X315 1 2 ICV_3 $T=161120 216000 0 0 $X=160830 $Y=215765
X316 1 2 ICV_3 $T=199200 200320 0 0 $X=198910 $Y=200085
X317 1 2 ICV_3 $T=199200 208160 0 0 $X=198910 $Y=207925
X318 1 2 ICV_3 $T=199200 223840 0 0 $X=198910 $Y=223605
X319 1 2 ICV_3 $T=210400 216000 1 0 $X=210110 $Y=211790
X320 1 2 ICV_3 $T=215440 223840 0 0 $X=215150 $Y=223605
X321 1 2 ICV_3 $T=216560 200320 0 0 $X=216270 $Y=200085
X322 1 2 ICV_3 $T=218800 208160 0 0 $X=218510 $Y=207925
X323 1 2 ICV_3 $T=225520 223840 1 0 $X=225230 $Y=219630
X324 1 2 ICV_3 $T=233360 231680 1 0 $X=233070 $Y=227470
X325 1 2 ICV_3 $T=241200 216000 1 0 $X=240910 $Y=211790
X326 1 2 ICV_3 $T=260800 216000 0 0 $X=260510 $Y=215765
X327 1 2 ICV_3 $T=277040 223840 1 0 $X=276750 $Y=219630
X328 1 2 ICV_3 $T=283200 208160 1 0 $X=282910 $Y=203950
X329 1 2 ICV_3 $T=283200 231680 1 0 $X=282910 $Y=227470
X330 1 2 ICV_3 $T=287120 223840 0 0 $X=286830 $Y=223605
X331 1 2 ICV_3 $T=309520 208160 0 0 $X=309230 $Y=207925
X332 1 2 ICV_3 $T=312880 231680 1 0 $X=312590 $Y=227470
X333 1 2 ICV_3 $T=318480 200320 0 0 $X=318190 $Y=200085
X334 1 2 ICV_3 $T=325200 231680 1 0 $X=324910 $Y=227470
X335 1 2 ICV_3 $T=329120 216000 1 0 $X=328830 $Y=211790
X336 1 2 ICV_3 $T=333600 208160 1 0 $X=333310 $Y=203950
X337 1 2 ICV_3 $T=347600 208160 1 0 $X=347310 $Y=203950
X338 1 2 ICV_3 $T=355440 216000 0 0 $X=355150 $Y=215765
X339 1 2 ICV_3 $T=358800 223840 0 0 $X=358510 $Y=223605
X340 1 2 ICV_3 $T=361600 223840 1 0 $X=361310 $Y=219630
X341 1 2 ICV_3 $T=371120 223840 0 0 $X=370830 $Y=223605
X342 1 2 ICV_3 $T=409200 200320 0 0 $X=408910 $Y=200085
X343 1 2 ICV_3 $T=409200 208160 1 0 $X=408910 $Y=203950
X344 1 2 ICV_3 $T=426560 208160 1 0 $X=426270 $Y=203950
X345 1 2 ICV_3 $T=433280 208160 0 0 $X=432990 $Y=207925
X346 1 2 ICV_3 $T=439440 216000 1 0 $X=439150 $Y=211790
X347 1 2 ICV_3 $T=441680 231680 1 0 $X=441390 $Y=227470
X348 1 2 ICV_3 $T=446160 208160 0 0 $X=445870 $Y=207925
X349 1 2 ICV_3 $T=451200 208160 0 0 $X=450910 $Y=207925
X350 1 2 ICV_3 $T=451200 223840 0 0 $X=450910 $Y=223605
X351 1 2 ICV_3 $T=455120 208160 1 0 $X=454830 $Y=203950
X352 1 2 ICV_3 $T=464640 208160 1 0 $X=464350 $Y=203950
X353 1 2 ICV_3 $T=465200 216000 1 0 $X=464910 $Y=211790
X354 1 2 DCAP8BWP7T $T=23920 216000 1 0 $X=23630 $Y=211790
X355 1 2 DCAP8BWP7T $T=29520 208160 0 0 $X=29230 $Y=207925
X356 1 2 DCAP8BWP7T $T=29520 231680 1 0 $X=29230 $Y=227470
X357 1 2 DCAP8BWP7T $T=59760 200320 0 0 $X=59470 $Y=200085
X358 1 2 DCAP8BWP7T $T=63680 223840 0 0 $X=63390 $Y=223605
X359 1 2 DCAP8BWP7T $T=84400 208160 1 0 $X=84110 $Y=203950
X360 1 2 DCAP8BWP7T $T=85520 216000 0 0 $X=85230 $Y=215765
X361 1 2 DCAP8BWP7T $T=101200 208160 1 0 $X=100910 $Y=203950
X362 1 2 DCAP8BWP7T $T=113520 208160 1 0 $X=113230 $Y=203950
X363 1 2 DCAP8BWP7T $T=125280 208160 1 0 $X=124990 $Y=203950
X364 1 2 DCAP8BWP7T $T=135360 208160 0 0 $X=135070 $Y=207925
X365 1 2 DCAP8BWP7T $T=142080 200320 0 0 $X=141790 $Y=200085
X366 1 2 DCAP8BWP7T $T=147120 216000 0 0 $X=146830 $Y=215765
X367 1 2 DCAP8BWP7T $T=152160 208160 0 0 $X=151870 $Y=207925
X368 1 2 DCAP8BWP7T $T=153280 200320 0 0 $X=152990 $Y=200085
X369 1 2 DCAP8BWP7T $T=153280 223840 1 0 $X=152990 $Y=219630
X370 1 2 DCAP8BWP7T $T=153840 208160 1 0 $X=153550 $Y=203950
X371 1 2 DCAP8BWP7T $T=153840 216000 0 0 $X=153550 $Y=215765
X372 1 2 DCAP8BWP7T $T=155520 223840 0 0 $X=155230 $Y=223605
X373 1 2 DCAP8BWP7T $T=184080 231680 1 0 $X=183790 $Y=227470
X374 1 2 DCAP8BWP7T $T=188000 216000 1 0 $X=187710 $Y=211790
X375 1 2 DCAP8BWP7T $T=196400 216000 0 0 $X=196110 $Y=215765
X376 1 2 DCAP8BWP7T $T=212080 200320 0 0 $X=211790 $Y=200085
X377 1 2 DCAP8BWP7T $T=212080 216000 0 0 $X=211790 $Y=215765
X378 1 2 DCAP8BWP7T $T=221600 200320 0 0 $X=221310 $Y=200085
X379 1 2 DCAP8BWP7T $T=225520 208160 1 0 $X=225230 $Y=203950
X380 1 2 DCAP8BWP7T $T=227200 231680 1 0 $X=226910 $Y=227470
X381 1 2 DCAP8BWP7T $T=239520 200320 0 0 $X=239230 $Y=200085
X382 1 2 DCAP8BWP7T $T=239520 208160 0 0 $X=239230 $Y=207925
X383 1 2 DCAP8BWP7T $T=239520 231680 1 0 $X=239230 $Y=227470
X384 1 2 DCAP8BWP7T $T=257440 208160 1 0 $X=257150 $Y=203950
X385 1 2 DCAP8BWP7T $T=266960 216000 0 0 $X=266670 $Y=215765
X386 1 2 DCAP8BWP7T $T=272560 223840 1 0 $X=272270 $Y=219630
X387 1 2 DCAP8BWP7T $T=277600 208160 0 0 $X=277310 $Y=207925
X388 1 2 DCAP8BWP7T $T=278720 208160 1 0 $X=278430 $Y=203950
X389 1 2 DCAP8BWP7T $T=280960 223840 0 0 $X=280670 $Y=223605
X390 1 2 DCAP8BWP7T $T=294400 216000 0 0 $X=294110 $Y=215765
X391 1 2 DCAP8BWP7T $T=297200 208160 1 0 $X=296910 $Y=203950
X392 1 2 DCAP8BWP7T $T=298880 223840 0 0 $X=298590 $Y=223605
X393 1 2 DCAP8BWP7T $T=301120 216000 1 0 $X=300830 $Y=211790
X394 1 2 DCAP8BWP7T $T=306720 208160 1 0 $X=306430 $Y=203950
X395 1 2 DCAP8BWP7T $T=311760 216000 1 0 $X=311470 $Y=211790
X396 1 2 DCAP8BWP7T $T=314000 200320 0 0 $X=313710 $Y=200085
X397 1 2 DCAP8BWP7T $T=317360 223840 0 0 $X=317070 $Y=223605
X398 1 2 DCAP8BWP7T $T=322960 216000 0 0 $X=322670 $Y=215765
X399 1 2 DCAP8BWP7T $T=323520 200320 0 0 $X=323230 $Y=200085
X400 1 2 DCAP8BWP7T $T=340880 231680 1 0 $X=340590 $Y=227470
X401 1 2 DCAP8BWP7T $T=343120 208160 1 0 $X=342830 $Y=203950
X402 1 2 DCAP8BWP7T $T=352640 216000 1 0 $X=352350 $Y=211790
X403 1 2 DCAP8BWP7T $T=356560 208160 1 0 $X=356270 $Y=203950
X404 1 2 DCAP8BWP7T $T=361600 216000 0 0 $X=361310 $Y=215765
X405 1 2 DCAP8BWP7T $T=362160 208160 0 0 $X=361870 $Y=207925
X406 1 2 DCAP8BWP7T $T=364400 223840 0 0 $X=364110 $Y=223605
X407 1 2 DCAP8BWP7T $T=364960 216000 1 0 $X=364670 $Y=211790
X408 1 2 DCAP8BWP7T $T=365520 208160 1 0 $X=365230 $Y=203950
X409 1 2 DCAP8BWP7T $T=376720 216000 1 0 $X=376430 $Y=211790
X410 1 2 DCAP8BWP7T $T=380080 223840 1 0 $X=379790 $Y=219630
X411 1 2 DCAP8BWP7T $T=381760 208160 0 0 $X=381470 $Y=207925
X412 1 2 DCAP8BWP7T $T=386240 223840 0 0 $X=385950 $Y=223605
X413 1 2 DCAP8BWP7T $T=387920 200320 0 0 $X=387630 $Y=200085
X414 1 2 DCAP8BWP7T $T=388480 223840 1 0 $X=388190 $Y=219630
X415 1 2 DCAP8BWP7T $T=393520 231680 1 0 $X=393230 $Y=227470
X416 1 2 DCAP8BWP7T $T=395200 223840 0 0 $X=394910 $Y=223605
X417 1 2 DCAP8BWP7T $T=402480 208160 0 0 $X=402190 $Y=207925
X418 1 2 DCAP8BWP7T $T=403600 216000 1 0 $X=403310 $Y=211790
X419 1 2 DCAP8BWP7T $T=407520 216000 0 0 $X=407230 $Y=215765
X420 1 2 DCAP8BWP7T $T=420400 216000 0 0 $X=420110 $Y=215765
X421 1 2 DCAP8BWP7T $T=423200 216000 1 0 $X=422910 $Y=211790
X422 1 2 DCAP8BWP7T $T=426560 200320 0 0 $X=426270 $Y=200085
X423 1 2 DCAP8BWP7T $T=427120 231680 1 0 $X=426830 $Y=227470
X424 1 2 DCAP8BWP7T $T=428800 208160 0 0 $X=428510 $Y=207925
X425 1 2 DCAP8BWP7T $T=429920 216000 0 0 $X=429630 $Y=215765
X426 1 2 DCAP8BWP7T $T=434400 208160 1 0 $X=434110 $Y=203950
X427 1 2 DCAP8BWP7T $T=434960 216000 1 0 $X=434670 $Y=211790
X428 1 2 DCAP8BWP7T $T=438880 208160 0 0 $X=438590 $Y=207925
X429 1 2 DCAP8BWP7T $T=445600 216000 1 0 $X=445310 $Y=211790
X430 1 2 DCAP8BWP7T $T=446160 231680 1 0 $X=445870 $Y=227470
X431 1 2 DCAP8BWP7T $T=447840 208160 1 0 $X=447550 $Y=203950
X432 1 2 DCAP8BWP7T $T=448400 200320 0 0 $X=448110 $Y=200085
X433 2 1 DCAPBWP7T $T=21120 200320 0 0 $X=20830 $Y=200085
X434 2 1 DCAPBWP7T $T=21120 208160 0 0 $X=20830 $Y=207925
X435 2 1 DCAPBWP7T $T=25600 208160 1 0 $X=25310 $Y=203950
X436 2 1 DCAPBWP7T $T=27840 216000 0 0 $X=27550 $Y=215765
X437 2 1 DCAPBWP7T $T=48000 216000 0 0 $X=47710 $Y=215765
X438 2 1 DCAPBWP7T $T=51920 208160 1 0 $X=51630 $Y=203950
X439 2 1 DCAPBWP7T $T=68160 223840 0 0 $X=67870 $Y=223605
X440 2 1 DCAPBWP7T $T=79360 208160 1 0 $X=79070 $Y=203950
X441 2 1 DCAPBWP7T $T=82720 208160 0 0 $X=82430 $Y=207925
X442 2 1 DCAPBWP7T $T=129760 200320 0 0 $X=129470 $Y=200085
X443 2 1 DCAPBWP7T $T=149360 200320 0 0 $X=149070 $Y=200085
X444 2 1 DCAPBWP7T $T=158320 208160 1 0 $X=158030 $Y=203950
X445 2 1 DCAPBWP7T $T=158320 216000 0 0 $X=158030 $Y=215765
X446 2 1 DCAPBWP7T $T=168400 208160 1 0 $X=168110 $Y=203950
X447 2 1 DCAPBWP7T $T=179040 200320 0 0 $X=178750 $Y=200085
X448 2 1 DCAPBWP7T $T=180720 216000 1 0 $X=180430 $Y=211790
X449 2 1 DCAPBWP7T $T=195840 208160 1 0 $X=195550 $Y=203950
X450 2 1 DCAPBWP7T $T=205360 231680 1 0 $X=205070 $Y=227470
X451 2 1 DCAPBWP7T $T=219360 231680 1 0 $X=219070 $Y=227470
X452 2 1 DCAPBWP7T $T=232800 223840 0 0 $X=232510 $Y=223605
X453 2 1 DCAPBWP7T $T=257440 231680 1 0 $X=257150 $Y=227470
X454 2 1 DCAPBWP7T $T=271440 216000 0 0 $X=271150 $Y=215765
X455 2 1 DCAPBWP7T $T=305600 216000 1 0 $X=305310 $Y=211790
X456 2 1 DCAPBWP7T $T=306160 208160 0 0 $X=305870 $Y=207925
X457 2 1 DCAPBWP7T $T=326320 208160 0 0 $X=326030 $Y=207925
X458 2 1 DCAPBWP7T $T=333600 200320 0 0 $X=333310 $Y=200085
X459 2 1 DCAPBWP7T $T=333600 208160 0 0 $X=333310 $Y=207925
X460 2 1 DCAPBWP7T $T=347600 216000 1 0 $X=347310 $Y=211790
X461 2 1 DCAPBWP7T $T=357120 216000 1 0 $X=356830 $Y=211790
X462 2 1 DCAPBWP7T $T=368320 231680 1 0 $X=368030 $Y=227470
X463 2 1 DCAPBWP7T $T=379520 200320 0 0 $X=379230 $Y=200085
X464 2 1 DCAPBWP7T $T=381200 216000 1 0 $X=380910 $Y=211790
X465 2 1 DCAPBWP7T $T=386240 208160 0 0 $X=385950 $Y=207925
X466 2 1 DCAPBWP7T $T=410320 223840 1 0 $X=410030 $Y=219630
X467 2 1 DCAPBWP7T $T=422080 231680 1 0 $X=421790 $Y=227470
X468 2 1 DCAPBWP7T $T=447280 216000 0 0 $X=446990 $Y=215765
X469 2 1 DCAPBWP7T $T=452320 208160 1 0 $X=452030 $Y=203950
X470 2 1 DCAPBWP7T $T=464080 200320 0 0 $X=463790 $Y=200085
X471 2 1 DCAPBWP7T $T=469120 223840 0 0 $X=468830 $Y=223605
X472 278 279 269 283 254 233 1 2 289 AO222D0BWP7T $T=234480 223840 1 0 $X=234190 $Y=219630
X473 279 278 291 294 295 233 1 2 297 AO222D0BWP7T $T=247920 216000 0 0 $X=247630 $Y=215765
X474 279 278 292 293 296 233 1 2 300 AO222D0BWP7T $T=248480 208160 0 0 $X=248190 $Y=207925
X475 278 279 292 301 299 233 1 2 290 AO222D0BWP7T $T=257440 231680 0 180 $X=250990 $Y=227470
X476 394 423 445 333 296 329 1 2 946 AO222D0BWP7T $T=364960 216000 0 180 $X=358510 $Y=211790
X477 476 469 467 465 464 423 1 2 950 AO222D0BWP7T $T=389040 216000 0 180 $X=382590 $Y=211790
X478 476 469 478 364 479 423 1 2 482 AO222D0BWP7T $T=394080 200320 0 0 $X=393790 $Y=200085
X479 476 469 956 467 466 423 1 2 955 AO222D0BWP7T $T=401360 223840 0 180 $X=394910 $Y=219630
X480 476 469 480 484 485 423 1 2 954 AO222D0BWP7T $T=397440 216000 1 0 $X=397150 $Y=211790
X481 518 1 517 515 514 2 962 513 OAI221D1BWP7T $T=437760 223840 1 180 $X=432430 $Y=223605
X482 359 278 363 279 368 233 1 2 372 AO222D1BWP7T $T=292720 231680 1 0 $X=292430 $Y=227470
X483 424 423 333 925 419 329 1 2 414 AO222D1BWP7T $T=342000 200320 1 180 $X=334990 $Y=200085
X484 425 423 333 396 421 329 1 2 417 AO222D1BWP7T $T=343120 208160 0 180 $X=336110 $Y=203950
X485 450 423 333 447 444 329 1 2 439 AO222D1BWP7T $T=366640 200320 1 180 $X=359630 $Y=200085
X486 1 2 ICV_4 $T=30080 223840 0 0 $X=29790 $Y=223605
X487 1 2 ICV_4 $T=35120 208160 1 0 $X=34830 $Y=203950
X488 1 2 ICV_4 $T=39600 200320 0 0 $X=39310 $Y=200085
X489 1 2 ICV_4 $T=48000 223840 1 0 $X=47710 $Y=219630
X490 1 2 ICV_4 $T=58640 231680 1 0 $X=58350 $Y=227470
X491 1 2 ICV_4 $T=72080 216000 1 0 $X=71790 $Y=211790
X492 1 2 ICV_4 $T=86640 231680 1 0 $X=86350 $Y=227470
X493 1 2 ICV_4 $T=93360 231680 1 0 $X=93070 $Y=227470
X494 1 2 ICV_4 $T=145440 216000 1 0 $X=145150 $Y=211790
X495 1 2 ICV_4 $T=156080 216000 1 0 $X=155790 $Y=211790
X496 1 2 ICV_4 $T=161120 200320 0 0 $X=160830 $Y=200085
X497 1 2 ICV_4 $T=161120 208160 0 0 $X=160830 $Y=207925
X498 1 2 ICV_4 $T=207600 223840 1 0 $X=207310 $Y=219630
X499 1 2 ICV_4 $T=245120 223840 0 0 $X=244830 $Y=223605
X500 1 2 ICV_4 $T=249600 223840 1 0 $X=249310 $Y=219630
X501 1 2 ICV_4 $T=282080 208160 0 0 $X=281790 $Y=207925
X502 1 2 ICV_4 $T=287120 216000 1 0 $X=286830 $Y=211790
X503 1 2 ICV_4 $T=324080 208160 1 0 $X=323790 $Y=203950
X504 1 2 ICV_4 $T=324080 223840 0 0 $X=323790 $Y=223605
X505 1 2 ICV_4 $T=366080 216000 0 0 $X=365790 $Y=215765
X506 1 2 ICV_4 $T=371120 216000 1 0 $X=370830 $Y=211790
X507 1 2 ICV_4 $T=399680 223840 0 0 $X=399390 $Y=223605
X508 1 2 ICV_4 $T=408080 216000 1 0 $X=407790 $Y=211790
X509 1 2 ICV_4 $T=413120 208160 1 0 $X=412830 $Y=203950
X510 1 2 ICV_4 $T=450080 216000 1 0 $X=449790 $Y=211790
X511 1 2 ICV_4 $T=455120 223840 0 0 $X=454830 $Y=223605
X512 1 2 ICV_4 $T=459600 208160 0 0 $X=459310 $Y=207925
X513 1 2 ICV_4 $T=466880 208160 0 0 $X=466590 $Y=207925
X514 214 212 208 2 1 198 DFCNQD1BWP7T $T=182960 223840 1 180 $X=170350 $Y=223605
X515 214 876 208 2 1 201 DFCNQD1BWP7T $T=184080 231680 0 180 $X=171470 $Y=227470
X516 214 889 208 2 1 246 DFCNQD1BWP7T $T=219360 231680 0 180 $X=206750 $Y=227470
X517 441 946 435 2 1 892 DFCNQD1BWP7T $T=362160 208160 1 180 $X=349550 $Y=207925
X700 1 2 ICV_9 $T=34000 200320 0 0 $X=33710 $Y=200085
X701 1 2 ICV_9 $T=34000 223840 1 0 $X=33710 $Y=219630
X702 1 2 ICV_9 $T=34000 223840 0 0 $X=33710 $Y=223605
X703 1 2 ICV_9 $T=34000 231680 1 0 $X=33710 $Y=227470
X704 1 2 ICV_9 $T=118000 216000 1 0 $X=117710 $Y=211790
X705 1 2 ICV_9 $T=118000 223840 1 0 $X=117710 $Y=219630
X706 1 2 ICV_9 $T=118000 231680 1 0 $X=117710 $Y=227470
X707 1 2 ICV_9 $T=160000 223840 1 0 $X=159710 $Y=219630
X708 1 2 ICV_9 $T=202000 208160 1 0 $X=201710 $Y=203950
X709 1 2 ICV_9 $T=202000 223840 1 0 $X=201710 $Y=219630
X710 1 2 ICV_9 $T=244000 223840 1 0 $X=243710 $Y=219630
X711 1 2 ICV_9 $T=286000 208160 1 0 $X=285710 $Y=203950
X712 1 2 ICV_9 $T=286000 208160 0 0 $X=285710 $Y=207925
X713 1 2 ICV_9 $T=286000 231680 1 0 $X=285710 $Y=227470
X714 1 2 ICV_9 $T=328000 200320 0 0 $X=327710 $Y=200085
X715 1 2 ICV_9 $T=328000 208160 1 0 $X=327710 $Y=203950
X716 1 2 ICV_9 $T=328000 208160 0 0 $X=327710 $Y=207925
X717 1 2 ICV_9 $T=328000 216000 0 0 $X=327710 $Y=215765
X718 1 2 ICV_9 $T=328000 223840 0 0 $X=327710 $Y=223605
X719 1 2 ICV_9 $T=328000 231680 1 0 $X=327710 $Y=227470
X720 1 2 ICV_9 $T=370000 200320 0 0 $X=369710 $Y=200085
X721 1 2 ICV_9 $T=370000 216000 0 0 $X=369710 $Y=215765
X722 1 2 ICV_9 $T=412000 200320 0 0 $X=411710 $Y=200085
X723 1 2 ICV_9 $T=412000 216000 1 0 $X=411710 $Y=211790
X724 1 2 ICV_9 $T=454000 208160 0 0 $X=453710 $Y=207925
X725 1 2 ICV_9 $T=454000 231680 1 0 $X=453710 $Y=227470
X726 1 2 ICV_13 $T=30640 200320 0 0 $X=30350 $Y=200085
X727 1 2 ICV_13 $T=30640 208160 1 0 $X=30350 $Y=203950
X728 1 2 ICV_13 $T=35120 208160 0 0 $X=34830 $Y=207925
X729 1 2 ICV_13 $T=35120 216000 0 0 $X=34830 $Y=215765
X730 1 2 ICV_13 $T=39600 231680 1 0 $X=39310 $Y=227470
X731 1 2 ICV_13 $T=42960 208160 1 0 $X=42670 $Y=203950
X732 1 2 ICV_13 $T=47440 200320 0 0 $X=47150 $Y=200085
X733 1 2 ICV_13 $T=56960 223840 0 0 $X=56670 $Y=223605
X734 1 2 ICV_13 $T=58640 208160 1 0 $X=58350 $Y=203950
X735 1 2 ICV_13 $T=86080 200320 0 0 $X=85790 $Y=200085
X736 1 2 ICV_13 $T=105680 208160 1 0 $X=105390 $Y=203950
X737 1 2 ICV_13 $T=114640 223840 0 0 $X=114350 $Y=223605
X738 1 2 ICV_13 $T=119120 216000 0 0 $X=118830 $Y=215765
X739 1 2 ICV_13 $T=123600 231680 1 0 $X=123310 $Y=227470
X740 1 2 ICV_13 $T=156640 208160 0 0 $X=156350 $Y=207925
X741 1 2 ICV_13 $T=161120 208160 1 0 $X=160830 $Y=203950
X742 1 2 ICV_13 $T=161120 223840 0 0 $X=160830 $Y=223605
X743 1 2 ICV_13 $T=192480 216000 1 0 $X=192190 $Y=211790
X744 1 2 ICV_13 $T=203120 208160 0 0 $X=202830 $Y=207925
X745 1 2 ICV_13 $T=203120 223840 0 0 $X=202830 $Y=223605
X746 1 2 ICV_13 $T=226640 208160 0 0 $X=226350 $Y=207925
X747 1 2 ICV_13 $T=245120 208160 0 0 $X=244830 $Y=207925
X748 1 2 ICV_13 $T=272000 208160 0 0 $X=271710 $Y=207925
X749 1 2 ICV_13 $T=298880 216000 0 0 $X=298590 $Y=215765
X750 1 2 ICV_13 $T=301120 223840 1 0 $X=300830 $Y=219630
X751 1 2 ICV_13 $T=306160 231680 1 0 $X=305870 $Y=227470
X752 1 2 ICV_13 $T=316800 216000 0 0 $X=316510 $Y=215765
X753 1 2 ICV_13 $T=366640 208160 0 0 $X=366350 $Y=207925
X754 1 2 ICV_13 $T=371120 208160 0 0 $X=370830 $Y=207925
X755 1 2 ICV_13 $T=408640 223840 0 0 $X=408350 $Y=223605
X756 1 2 ICV_13 $T=413120 223840 0 0 $X=412830 $Y=223605
X757 1 2 ICV_13 $T=429360 223840 0 0 $X=429070 $Y=223605
X758 1 2 ICV_13 $T=431600 231680 1 0 $X=431310 $Y=227470
X759 1 2 ICV_13 $T=450640 216000 0 0 $X=450350 $Y=215765
X760 1 2 ICV_13 $T=450640 231680 1 0 $X=450350 $Y=227470
X761 1 2 ICV_13 $T=455120 216000 1 0 $X=454830 $Y=211790
X762 387 390 2 390 927 387 1 MAOI22D1BWP7T $T=311760 216000 0 180 $X=306990 $Y=211790
X763 351 233 1 347 346 2 IOA21D0BWP7T $T=283200 231680 0 180 $X=279550 $Y=227470
X764 505 344 1 960 502 2 IOA21D0BWP7T $T=427120 231680 0 180 $X=423470 $Y=227470
X765 4 1 2 772 INVD1BWP7T $T=22240 216000 1 0 $X=21950 $Y=211790
X766 58 1 2 57 INVD1BWP7T $T=58640 208160 0 180 $X=56670 $Y=203950
X767 68 1 2 55 INVD1BWP7T $T=66480 216000 0 0 $X=66190 $Y=215765
X768 89 1 2 792 INVD1BWP7T $T=86640 231680 0 180 $X=84670 $Y=227470
X769 90 1 2 799 INVD1BWP7T $T=91680 208160 0 0 $X=91390 $Y=207925
X770 114 1 2 128 INVD1BWP7T $T=130320 223840 1 180 $X=128350 $Y=223605
X771 130 1 2 143 INVD1BWP7T $T=138160 216000 0 180 $X=136190 $Y=211790
X772 845 1 2 146 INVD1BWP7T $T=138720 223840 0 0 $X=138430 $Y=223605
X773 867 1 2 200 INVD1BWP7T $T=170080 231680 1 0 $X=169790 $Y=227470
X774 172 1 2 298 INVD1BWP7T $T=255200 223840 0 180 $X=253230 $Y=219630
X775 362 1 2 917 INVD1BWP7T $T=294400 223840 1 180 $X=292430 $Y=223605
X776 391 1 2 393 INVD1BWP7T $T=312320 200320 0 0 $X=312030 $Y=200085
X777 392 1 2 397 INVD1BWP7T $T=312320 208160 0 0 $X=312030 $Y=207925
X778 396 1 2 398 INVD1BWP7T $T=319600 208160 1 180 $X=317630 $Y=207925
X779 937 1 2 412 INVD1BWP7T $T=335840 223840 1 180 $X=333870 $Y=223605
X780 550 544 1 2 BUFFD2BWP7T $T=468000 231680 0 180 $X=464350 $Y=227470
X781 561 549 1 2 BUFFD2BWP7T $T=470800 208160 0 180 $X=467150 $Y=203950
X782 1 2 DCAP16BWP7T $T=21120 223840 0 0 $X=20830 $Y=223605
X783 1 2 DCAP16BWP7T $T=55280 216000 1 0 $X=54990 $Y=211790
X784 1 2 DCAP16BWP7T $T=161120 231680 1 0 $X=160830 $Y=227470
X785 1 2 DCAP16BWP7T $T=203120 216000 0 0 $X=202830 $Y=215765
X786 1 2 DCAP16BWP7T $T=245120 208160 1 0 $X=244830 $Y=203950
X787 1 2 DCAP16BWP7T $T=340320 208160 0 0 $X=340030 $Y=207925
X788 1 2 DCAP16BWP7T $T=389600 216000 0 0 $X=389310 $Y=215765
X789 1 2 DCAP16BWP7T $T=400240 200320 0 0 $X=399950 $Y=200085
X790 1 2 DCAP16BWP7T $T=401360 223840 1 0 $X=401070 $Y=219630
X791 1 2 DCAP16BWP7T $T=420400 223840 0 0 $X=420110 $Y=223605
X792 1 2 DCAP16BWP7T $T=429360 223840 1 0 $X=429070 $Y=219630
X793 1 2 DCAP16BWP7T $T=433280 200320 0 0 $X=432990 $Y=200085
X794 1 2 DCAP16BWP7T $T=437760 223840 0 0 $X=437470 $Y=223605
X795 1 2 DCAP16BWP7T $T=445040 223840 1 0 $X=444750 $Y=219630
X796 1 2 DCAP16BWP7T $T=455120 200320 0 0 $X=454830 $Y=200085
X797 800 1 2 789 CKND1BWP7T $T=71520 223840 1 180 $X=69550 $Y=223605
X798 819 1 2 827 CKND1BWP7T $T=102880 223840 1 0 $X=102590 $Y=219630
X799 131 1 2 843 CKND1BWP7T $T=121920 208160 0 0 $X=121630 $Y=207925
X800 183 1 2 862 CKND1BWP7T $T=153840 216000 1 180 $X=151870 $Y=215765
X801 178 1 2 195 CKND1BWP7T $T=168960 208160 0 0 $X=168670 $Y=207925
X802 313 1 2 331 CKND1BWP7T $T=272000 231680 1 0 $X=271710 $Y=227470
X803 389 1 2 376 CKND1BWP7T $T=309520 208160 1 180 $X=307550 $Y=207925
X804 860 1 2 418 CKND1BWP7T $T=332480 223840 1 0 $X=332190 $Y=219630
X805 866 1 2 216 BUFFD3BWP7T $T=186880 223840 1 180 $X=182670 $Y=223605
X806 878 1 2 260 BUFFD3BWP7T $T=213200 216000 1 0 $X=212910 $Y=211790
X807 271 873 2 895 1 273 899 AOI22D1BWP7T $T=226640 223840 0 0 $X=226350 $Y=223605
X808 277 897 2 276 1 893 898 AOI22D1BWP7T $T=233920 208160 1 180 $X=229710 $Y=207925
X809 329 299 2 333 1 338 334 AOI22D1BWP7T $T=279840 231680 0 180 $X=275630 $Y=227470
X810 329 341 2 333 1 348 349 AOI22D1BWP7T $T=278160 200320 0 0 $X=277870 $Y=200085
X811 440 437 2 443 1 446 947 AOI22D1BWP7T $T=359920 231680 1 0 $X=359630 $Y=227470
X812 329 434 2 333 1 448 944 AOI22D1BWP7T $T=361600 208160 1 0 $X=361310 $Y=203950
X813 475 473 2 472 1 470 952 AOI22D1BWP7T $T=393520 231680 0 180 $X=389310 $Y=227470
X814 477 473 2 474 1 470 471 AOI22D1BWP7T $T=395200 223840 1 180 $X=390990 $Y=223605
X815 191 184 2 863 188 1 OAI21D1BWP7T $T=168400 200320 1 180 $X=164750 $Y=200085
X816 256 878 2 888 253 1 OAI21D1BWP7T $T=214880 223840 0 180 $X=211230 $Y=219630
X817 315 260 2 914 317 1 OAI21D1BWP7T $T=263600 216000 0 0 $X=263310 $Y=215765
X818 394 930 2 931 928 1 OAI21D1BWP7T $T=313440 216000 0 0 $X=313150 $Y=215765
X819 244 233 1 2 BUFFD8BWP7T $T=206480 223840 0 0 $X=206190 $Y=223605
X820 868 2 190 186 1 NR2D4BWP7T $T=174000 216000 1 180 $X=166990 $Y=215765
X821 9 5 2 1 INVD2BWP7T $T=23360 231680 0 180 $X=20830 $Y=227470
X822 182 173 2 1 INVD2BWP7T $T=153280 200320 1 180 $X=150750 $Y=200085
X823 210 176 2 1 INVD2BWP7T $T=176800 216000 0 180 $X=174270 $Y=211790
X824 261 383 2 1 INVD2BWP7T $T=304480 208160 1 0 $X=304190 $Y=203950
X825 382 327 2 1 INVD2BWP7T $T=305040 223840 1 0 $X=304750 $Y=219630
X826 434 433 2 1 INVD2BWP7T $T=353200 200320 1 180 $X=350670 $Y=200085
X827 510 511 2 1 INVD2BWP7T $T=431040 200320 0 0 $X=430750 $Y=200085
X828 259 873 1 2 895 CKXOR2D1BWP7T $T=218240 223840 0 0 $X=217950 $Y=223605
X829 262 873 1 2 893 CKXOR2D1BWP7T $T=220480 223840 1 0 $X=220190 $Y=219630
X830 291 172 1 2 908 CKXOR2D1BWP7T $T=249040 223840 0 0 $X=248750 $Y=223605
X831 908 336 1 2 918 CKXOR2D1BWP7T $T=273120 216000 0 0 $X=272830 $Y=215765
X832 364 261 1 2 375 CKXOR2D1BWP7T $T=296080 223840 1 0 $X=295790 $Y=219630
X833 860 415 1 2 934 CKXOR2D1BWP7T $T=331920 216000 1 0 $X=331630 $Y=211790
X834 934 420 1 2 935 CKXOR2D1BWP7T $T=335280 208160 0 0 $X=334990 $Y=207925
X835 422 418 1 2 416 CKXOR2D1BWP7T $T=340880 231680 0 180 $X=335550 $Y=227470
X836 489 480 1 2 957 CKXOR2D1BWP7T $T=403600 223840 0 0 $X=403310 $Y=223605
X837 957 498 1 2 958 CKXOR2D1BWP7T $T=423200 216000 0 180 $X=417870 $Y=211790
X838 959 512 1 2 961 CKXOR2D1BWP7T $T=429360 208160 1 0 $X=429070 $Y=203950
X839 890 254 252 1 2 CKXOR2D2BWP7T $T=218800 208160 1 180 $X=212350 $Y=207925
X840 405 932 395 1 2 CKXOR2D2BWP7T $T=321280 223840 0 180 $X=314830 $Y=219630
X841 434 940 431 1 2 CKXOR2D2BWP7T $T=356560 208160 0 180 $X=350110 $Y=203950
X842 960 499 501 1 2 CKXOR2D2BWP7T $T=428800 208160 1 180 $X=422350 $Y=207925
X843 194 863 176 196 1 2 OAI21D0BWP7T $T=168400 200320 0 0 $X=168110 $Y=200085
X844 896 929 381 924 1 2 OAI21D0BWP7T $T=312880 231680 0 180 $X=309790 $Y=227470
X845 943 942 436 945 1 2 OAI21D0BWP7T $T=356000 223840 0 0 $X=355710 $Y=223605
X846 947 948 449 277 1 2 OAI21D0BWP7T $T=376160 223840 0 0 $X=375870 $Y=223605
X847 953 951 458 277 1 2 OAI21D0BWP7T $T=382320 223840 1 180 $X=379230 $Y=223605
X848 401 399 404 1 2 411 MUX2ND1BWP7T $T=316800 216000 1 0 $X=316510 $Y=211790
X849 893 256 1 2 897 XNR2D1BWP7T $T=220480 216000 1 0 $X=220190 $Y=211790
X850 269 266 1 2 894 XNR2D1BWP7T $T=226640 208160 1 180 $X=221310 $Y=207925
X851 270 272 1 2 275 XNR2D1BWP7T $T=226080 200320 0 0 $X=225790 $Y=200085
X852 275 903 1 2 901 XNR2D1BWP7T $T=234480 200320 0 0 $X=234190 $Y=200085
X853 280 904 1 2 905 XNR2D1BWP7T $T=234480 223840 0 0 $X=234190 $Y=223605
X854 313 309 1 2 177 XNR2D1BWP7T $T=263040 223840 1 180 $X=257710 $Y=223605
X855 495 891 1 2 959 XNR2D1BWP7T $T=417040 208160 1 0 $X=416750 $Y=203950
X856 503 904 2 1 CKND2BWP7T $T=434960 216000 0 180 $X=432430 $Y=211790
X857 365 1 2 356 CKND0BWP7T $T=293280 208160 0 180 $X=291310 $Y=203950
X858 367 1 2 903 CKND0BWP7T $T=297200 208160 0 180 $X=295230 $Y=203950
X859 493 1 2 488 CKND0BWP7T $T=408640 208160 1 180 $X=406670 $Y=207925
X860 490 488 492 490 488 2 1 IAO22D1BWP7T $T=409200 208160 0 180 $X=403870 $Y=203950
X861 195 2 197 882 182 880 1 AOI22D2BWP7T $T=181840 208160 0 0 $X=181550 $Y=207925
X862 277 2 901 284 275 276 1 AOI22D2BWP7T $T=230560 208160 1 0 $X=230270 $Y=203950
X863 298 2 906 307 303 172 1 AOI22D2BWP7T $T=252400 216000 1 0 $X=252110 $Y=211790
X864 302 2 298 312 172 310 1 AOI22D2BWP7T $T=254640 208160 0 0 $X=254350 $Y=207925
X865 329 2 328 330 335 333 1 AOI22D2BWP7T $T=272000 208160 1 0 $X=271710 $Y=203950
X866 329 2 361 352 354 333 1 AOI22D2BWP7T $T=296640 200320 1 180 $X=289630 $Y=200085
X867 329 2 254 914 423 936 1 AOI22D2BWP7T $T=347600 216000 0 180 $X=340590 $Y=211790
X868 427 2 329 888 423 426 1 AOI22D2BWP7T $T=347600 223840 0 180 $X=340590 $Y=219630
X869 329 2 466 460 461 333 1 AOI22D2BWP7T $T=387920 200320 1 180 $X=380910 $Y=200085
X870 956 2 481 494 487 483 1 AOI22D2BWP7T $T=398560 231680 1 0 $X=398270 $Y=227470
X871 486 2 481 491 487 484 1 AOI22D2BWP7T $T=400800 216000 0 0 $X=400510 $Y=215765
X872 329 2 496 920 503 333 1 AOI22D2BWP7T $T=419840 200320 0 0 $X=419550 $Y=200085
X873 895 274 900 902 1 2 MUX2ND0BWP7T $T=228320 223840 1 0 $X=228030 $Y=219630
X874 894 282 285 287 1 2 MUX2ND0BWP7T $T=235040 208160 0 0 $X=234750 $Y=207925
X875 817 147 146 139 36 2 1 AOI22D0BWP7T $T=133120 231680 0 180 $X=129470 $Y=227470
X876 184 883 220 228 884 2 1 AOI22D0BWP7T $T=190800 208160 0 0 $X=190510 $Y=207925
X877 905 286 280 277 276 2 1 AOI22D0BWP7T $T=239520 231680 0 180 $X=235870 $Y=227470
X878 163 1 2 164 CKBD0BWP7T $T=142080 231680 1 0 $X=141790 $Y=227470
X879 947 1 2 938 CKBD0BWP7T $T=361600 223840 0 180 $X=359070 $Y=219630
X880 197 195 202 869 2 1 206 AO211D1BWP7T $T=170640 208160 0 0 $X=170350 $Y=207925
X881 881 184 168 231 2 1 235 AO211D1BWP7T $T=191360 208160 1 0 $X=191070 $Y=203950
X882 6 2 771 3 1 NR2D1BWP7T $T=23360 208160 0 180 $X=20830 $Y=203950
X883 32 2 782 31 1 NR2D1BWP7T $T=42400 223840 0 180 $X=39870 $Y=219630
X884 37 2 784 61 1 NR2D1BWP7T $T=57520 200320 0 0 $X=57230 $Y=200085
X885 56 2 60 31 1 NR2D1BWP7T $T=60320 223840 0 180 $X=57790 $Y=219630
X886 52 2 797 75 1 NR2D1BWP7T $T=66480 208160 0 0 $X=66190 $Y=207925
X887 91 2 800 56 1 NR2D1BWP7T $T=88320 223840 0 180 $X=85790 $Y=219630
X888 103 2 801 105 1 NR2D1BWP7T $T=95600 200320 0 0 $X=95310 $Y=200085
X889 818 2 118 82 1 NR2D1BWP7T $T=107920 200320 0 0 $X=107630 $Y=200085
X890 838 2 129 55 1 NR2D1BWP7T $T=115200 200320 1 180 $X=112670 $Y=200085
X891 216 2 881 199 1 NR2D1BWP7T $T=184080 208160 1 0 $X=183790 $Y=203950
X892 211 2 884 881 1 NR2D1BWP7T $T=188560 208160 0 0 $X=188270 $Y=207925
X893 172 2 305 304 1 NR2D1BWP7T $T=258560 223840 0 180 $X=256030 $Y=219630
X894 860 2 407 409 1 NR2D1BWP7T $T=324080 223840 1 180 $X=321550 $Y=223605
X895 175 874 875 203 1 2 AOI21D0BWP7T $T=177920 216000 1 0 $X=177630 $Y=211790
X896 204 872 182 215 1 2 AOI21D0BWP7T $T=179040 208160 0 0 $X=178750 $Y=207925
X897 896 924 381 343 1 2 AOI21D0BWP7T $T=303360 231680 1 0 $X=303070 $Y=227470
X898 930 931 394 343 1 2 AOI21D0BWP7T $T=320160 216000 0 0 $X=319870 $Y=215765
X899 943 945 436 343 1 2 AOI21D0BWP7T $T=361600 223840 0 0 $X=361310 $Y=223605
X900 938 941 449 948 1 2 AOI21D0BWP7T $T=364400 223840 1 0 $X=364110 $Y=219630
X901 953 468 458 951 1 2 AOI21D0BWP7T $T=385680 223840 1 0 $X=385390 $Y=219630
X902 774 13 16 776 2 1 27 NR4D1BWP7T $T=23920 223840 1 0 $X=23630 $Y=219630
X903 824 101 789 815 2 1 40 NR4D1BWP7T $T=96160 223840 1 180 $X=90270 $Y=223605
X904 111 41 109 112 2 1 84 NR4D1BWP7T $T=98400 200320 0 0 $X=98110 $Y=200085
X905 832 84 115 48 2 1 820 NR4D1BWP7T $T=106800 231680 0 180 $X=100910 $Y=227470
X906 847 137 844 142 2 1 820 NR4D1BWP7T $T=123600 216000 1 0 $X=123310 $Y=211790
X907 89 59 90 798 2 1 814 OR4D1BWP7T $T=84960 216000 1 0 $X=84670 $Y=211790
X908 849 2 161 146 833 1 AOI21D2BWP7T $T=137040 216000 0 0 $X=136750 $Y=215765
X909 230 2 227 226 203 1 AOI21D2BWP7T $T=194160 200320 1 180 $X=188830 $Y=200085
X910 43 1 41 779 2 ND2D1BWP7T $T=51920 208160 0 180 $X=49390 $Y=203950
X911 29 1 82 69 2 ND2D1BWP7T $T=80480 208160 0 0 $X=80190 $Y=207925
X912 24 1 821 85 2 ND2D1BWP7T $T=89440 223840 1 0 $X=89150 $Y=219630
X913 72 1 820 102 2 ND2D1BWP7T $T=93360 216000 1 0 $X=93070 $Y=211790
X914 74 1 103 822 2 ND2D1BWP7T $T=98960 208160 0 180 $X=96430 $Y=203950
X915 92 1 811 74 2 ND2D1BWP7T $T=98960 208160 1 0 $X=98670 $Y=203950
X916 104 1 818 830 2 ND2D1BWP7T $T=104000 208160 0 0 $X=103710 $Y=207925
X917 166 1 130 857 2 ND2D1BWP7T $T=146560 231680 0 180 $X=144030 $Y=227470
X918 857 1 108 859 2 ND2D1BWP7T $T=146560 231680 1 0 $X=146270 $Y=227470
X919 177 1 845 166 2 ND2D1BWP7T $T=151040 231680 0 180 $X=148510 $Y=227470
X920 177 1 114 859 2 ND2D1BWP7T $T=154960 231680 0 180 $X=152430 $Y=227470
X921 837 1 846 832 2 849 108 OAI211D1BWP7T $T=124160 223840 1 0 $X=123870 $Y=219630
X922 205 1 870 207 2 869 184 OAI211D1BWP7T $T=173440 208160 1 0 $X=173150 $Y=203950
X923 868 1 864 190 2 871 210 OAI211D1BWP7T $T=174000 216000 0 0 $X=173710 $Y=215765
X924 224 1 227 884 2 229 178 OAI211D1BWP7T $T=189680 223840 1 0 $X=189390 $Y=219630
X925 224 1 227 884 2 232 178 OAI211D1BWP7T $T=191360 223840 0 0 $X=191070 $Y=223605
X926 247 1 248 203 2 249 207 OAI211D1BWP7T $T=210400 216000 0 180 $X=206750 $Y=211790
X927 265 1 267 894 2 890 268 OAI211D1BWP7T $T=222160 208160 1 0 $X=221870 $Y=203950
X928 928 1 386 385 2 922 345 OAI211D1BWP7T $T=308400 223840 1 180 $X=304750 $Y=223605
X929 942 1 429 428 2 937 345 OAI211D1BWP7T $T=350400 231680 0 180 $X=346750 $Y=227470
X930 463 1 462 952 2 457 345 OAI211D1BWP7T $T=384000 231680 0 180 $X=380350 $Y=227470
X931 773 2 27 781 789 1 790 NR4D2BWP7T $T=39600 223840 0 0 $X=39310 $Y=223605
X932 778 2 20 42 772 1 45 NR4D2BWP7T $T=42400 216000 1 0 $X=42110 $Y=211790
X933 178 2 189 194 1 NR2XD0BWP7T $T=166720 208160 0 0 $X=166430 $Y=207925
X934 190 2 196 880 1 NR2XD0BWP7T $T=181840 208160 1 0 $X=181550 $Y=203950
X935 7 1 10 771 8 773 2 ND4D1BWP7T $T=22800 200320 0 0 $X=22510 $Y=200085
X936 25 1 23 777 18 778 2 ND4D1BWP7T $T=30640 200320 1 180 $X=26430 $Y=200085
X937 780 1 24 23 30 781 2 ND4D1BWP7T $T=42960 208160 0 180 $X=38750 $Y=203950
X938 35 1 779 12 784 786 2 ND4D1BWP7T $T=43520 200320 0 0 $X=43230 $Y=200085
X939 38 1 785 774 30 36 2 ND4D1BWP7T $T=48000 223840 0 180 $X=43790 $Y=219630
X940 80 1 792 77 782 776 2 ND4D1BWP7T $T=71520 223840 0 180 $X=67310 $Y=219630
X941 68 1 24 792 799 812 2 ND4D1BWP7T $T=80480 223840 1 0 $X=80190 $Y=219630
X942 80 1 49 85 777 809 2 ND4D1BWP7T $T=85520 216000 1 180 $X=81310 $Y=215765
X943 117 827 837 120 128 1 2 OAI31D1BWP7T $T=108480 223840 1 0 $X=108190 $Y=219630
X944 119 827 841 813 128 1 2 OAI31D1BWP7T $T=110720 223840 0 0 $X=110430 $Y=223605
X945 791 138 846 786 143 1 2 OAI31D1BWP7T $T=125840 208160 0 0 $X=125550 $Y=207925
X946 66 155 152 848 128 1 2 OAI31D1BWP7T $T=136480 216000 0 180 $X=132270 $Y=211790
X947 24 1 797 50 2 802 ND3D0BWP7T $T=69280 216000 1 0 $X=68990 $Y=211790
X948 79 1 21 801 2 788 ND3D0BWP7T $T=72640 200320 1 180 $X=69550 $Y=200085
X949 68 1 810 88 2 813 ND3D0BWP7T $T=82720 223840 0 0 $X=82430 $Y=223605
X950 792 1 85 99 2 100 ND3D0BWP7T $T=90560 231680 1 0 $X=90270 $Y=227470
X951 92 1 106 782 2 825 ND3D0BWP7T $T=96720 216000 0 0 $X=96430 $Y=215765
X952 73 1 106 843 2 844 ND3D0BWP7T $T=123040 216000 0 0 $X=122750 $Y=215765
X953 213 1 190 176 2 877 ND3D0BWP7T $T=179040 208160 1 0 $X=178750 $Y=203950
X954 788 1 2 781 28 787 37 NR4D0BWP7T $T=49680 208160 0 180 $X=46030 $Y=203950
X955 811 1 2 84 57 810 42 NR4D0BWP7T $T=84400 208160 0 180 $X=80750 $Y=203950
X956 806 1 2 825 827 826 86 NR4D0BWP7T $T=99520 223840 1 0 $X=99230 $Y=219630
X957 816 1 2 110 825 828 112 NR4D0BWP7T $T=100080 216000 1 0 $X=99790 $Y=211790
X958 771 69 54 71 2 1 73 AN4D1BWP7T $T=64800 200320 0 0 $X=64510 $Y=200085
X959 800 98 72 85 2 1 819 AN4D1BWP7T $T=90560 216000 0 0 $X=90270 $Y=215765
X960 805 97 107 822 108 2 1 AOI31D1BWP7T $T=97280 231680 1 0 $X=96990 $Y=227470
X961 824 88 116 830 114 2 1 AOI31D1BWP7T $T=105120 223840 0 0 $X=104830 $Y=223605
X962 795 121 124 835 130 2 1 AOI31D1BWP7T $T=109600 231680 1 0 $X=109310 $Y=227470
X963 122 830 840 39 108 2 1 AOI31D1BWP7T $T=111280 216000 0 0 $X=110990 $Y=215765
X964 132 801 134 135 845 2 1 AOI31D1BWP7T $T=121920 200320 0 0 $X=121630 $Y=200085
X965 154 831 852 148 845 2 1 AOI31D1BWP7T $T=135360 200320 1 180 $X=131150 $Y=200085
X966 62 1 58 792 60 63 2 ND4D0BWP7T $T=63680 223840 1 180 $X=60030 $Y=223605
X967 58 1 72 24 74 798 2 ND4D0BWP7T $T=65920 216000 1 0 $X=65630 $Y=211790
X968 43 1 799 797 21 806 2 ND4D0BWP7T $T=69280 208160 1 0 $X=68990 $Y=203950
X969 76 1 78 800 803 804 2 ND4D0BWP7T $T=69280 216000 0 0 $X=68990 $Y=215765
X970 77 1 71 95 97 815 2 ND4D0BWP7T $T=89440 200320 0 0 $X=89150 $Y=200085
X971 92 1 807 94 803 817 2 ND4D0BWP7T $T=89440 216000 1 0 $X=89150 $Y=211790
X972 123 1 125 127 835 842 2 ND4D0BWP7T $T=111280 208160 0 0 $X=110990 $Y=207925
X973 133 1 96 831 843 136 2 ND4D0BWP7T $T=121920 208160 1 0 $X=121630 $Y=203950
X974 125 1 140 33 831 848 2 ND4D0BWP7T $T=126400 200320 0 0 $X=126110 $Y=200085
X975 838 1 811 821 831 2 NR3D1BWP7T $T=109040 208160 1 0 $X=108750 $Y=203950
X976 42 1 29 24 793 68 2 IND4D0BWP7T $T=59760 208160 0 0 $X=59470 $Y=207925
X977 791 1 97 104 823 72 2 IND4D0BWP7T $T=99520 216000 0 180 $X=95310 $Y=211790
X978 105 1 831 113 829 799 2 IND4D0BWP7T $T=107920 200320 1 180 $X=103710 $Y=200085
X979 31 1 46 49 791 51 2 IND4D1BWP7T $T=50800 200320 0 0 $X=50510 $Y=200085
X980 56 1 50 774 48 46 2 IND4D1BWP7T $T=56400 223840 0 180 $X=51630 $Y=219630
X981 811 1 87 83 808 8 2 IND4D1BWP7T $T=86080 200320 1 180 $X=81310 $Y=200085
X982 783 2 40 47 772 1 53 NR4D3BWP7T $T=42960 231680 1 0 $X=42670 $Y=227470
X983 64 793 66 47 2 1 796 OR4D0BWP7T $T=62000 216000 0 0 $X=61710 $Y=215765
X984 20 19 11 12 8 1 2 INR4D1BWP7T $T=29520 208160 1 180 $X=22510 $Y=207925
X985 55 37 59 785 62 1 2 INR4D1BWP7T $T=54720 216000 0 0 $X=54430 $Y=215765
X986 65 16 794 795 72 1 2 INR4D1BWP7T $T=62560 231680 1 0 $X=62270 $Y=227470
X987 110 821 126 839 80 1 2 INR4D1BWP7T $T=108480 216000 1 0 $X=108190 $Y=211790
X988 772 2 14 1 13 NR2XD1BWP7T $T=23920 216000 0 0 $X=23630 $Y=215765
X989 184 2 861 1 192 NR2XD1BWP7T $T=164480 208160 1 0 $X=164190 $Y=203950
X990 191 2 204 1 199 NR2XD1BWP7T $T=171200 200320 0 0 $X=170910 $Y=200085
X991 128 151 840 854 156 1 2 AO211D2BWP7T $T=132560 223840 1 0 $X=132270 $Y=219630
X992 143 162 852 856 165 1 2 AO211D2BWP7T $T=140400 216000 1 0 $X=140110 $Y=211790
X993 226 234 236 238 240 1 2 AO211D2BWP7T $T=194160 200320 0 0 $X=193870 $Y=200085
X994 875 1 878 216 2 194 879 OAI211D0BWP7T $T=184640 216000 1 180 $X=180990 $Y=215765
X995 886 1 882 210 2 207 887 OAI211D0BWP7T $T=195840 216000 1 0 $X=195550 $Y=211790
X996 929 1 402 933 2 345 932 OAI211D0BWP7T $T=317360 231680 1 0 $X=317070 $Y=227470
X997 342 1 939 432 2 268 940 OAI211D0BWP7T $T=349280 216000 1 0 $X=348990 $Y=211790
X998 880 1 194 878 2 CKND2D1BWP7T $T=184640 216000 0 180 $X=182110 $Y=211790
X999 865 1 864 187 193 173 2 OAI211D2BWP7T $T=170640 223840 1 180 $X=164190 $Y=223605
X1000 877 1 217 219 222 199 2 OAI211D2BWP7T $T=180720 200320 0 0 $X=180430 $Y=200085
X1001 886 1 882 207 243 210 2 OAI211D2BWP7T $T=193040 223840 1 0 $X=192750 $Y=219630
X1002 250 1 241 175 245 234 2 OAI211D2BWP7T $T=212080 200320 1 180 $X=205630 $Y=200085
X1003 247 1 248 207 251 203 2 OAI211D2BWP7T $T=206480 208160 0 0 $X=206190 $Y=207925
X1004 250 1 241 175 255 234 2 OAI211D2BWP7T $T=208720 208160 1 0 $X=208430 $Y=203950
X1005 898 1 899 902 288 281 2 OAI211D2BWP7T $T=230560 216000 1 0 $X=230270 $Y=211790
X1006 342 1 919 268 332 340 2 OAI211D2BWP7T $T=280960 216000 0 180 $X=274510 $Y=211790
X1007 204 203 874 871 1 2 867 AO211D0BWP7T $T=181280 216000 1 180 $X=177070 $Y=215765
X1008 221 213 215 883 1 2 885 AO211D0BWP7T $T=186880 208160 1 0 $X=186590 $Y=203950
X1009 233 2 230 886 204 221 1 AOI211D2BWP7T $T=196400 216000 1 180 $X=189950 $Y=215765
X1010 34 780 1 2 777 AN2D1BWP7T $T=41280 208160 1 180 $X=38190 $Y=207925
X1011 74 104 1 2 835 AN2D1BWP7T $T=106240 208160 0 0 $X=105950 $Y=207925
X1012 199 175 211 1 2 ND2D2BWP7T $T=175120 200320 0 0 $X=174830 $Y=200085
X1013 357 2 903 916 360 1 367 923 AOI221D1BWP7T $T=292160 208160 0 0 $X=291870 $Y=207925
X1014 357 2 376 377 379 1 925 926 AOI221D1BWP7T $T=300560 200320 0 0 $X=300270 $Y=200085
X1015 400 2 963 511 510 1 533 527 AOI221D1BWP7T $T=443360 200320 0 0 $X=443070 $Y=200085
X1016 802 1 2 81 59 807 NR3D0BWP7T $T=80480 216000 1 0 $X=80190 $Y=211790
X1017 344 350 1 353 919 2 AOI21D1BWP7T $T=279840 223840 1 0 $X=279550 $Y=219630
X1018 39 33 777 29 783 1 2 ND4D2BWP7T $T=45760 216000 1 180 $X=38190 $Y=215765
X1019 139 1 141 809 812 844 2 OAI31D2BWP7T $T=128640 223840 1 180 $X=121630 $Y=223605
X1020 26 1 24 21 2 19 ND3D1BWP7T $T=30640 208160 0 180 $X=26990 $Y=203950
X1021 203 1 191 199 2 868 ND3D1BWP7T $T=173440 208160 0 180 $X=169790 $Y=203950
X1022 868 1 209 870 2 873 ND3D1BWP7T $T=175120 208160 0 0 $X=174830 $Y=207925
X1023 941 2 430 938 1 939 276 AOI211D1BWP7T $T=350960 216000 1 180 $X=347310 $Y=215765
X1024 782 2 822 804 1 INR2D1BWP7T $T=99520 223840 0 180 $X=96430 $Y=219630
X1028 861 1 2 186 176 865 862 AOI211XD0BWP7T $T=163920 216000 0 0 $X=163630 $Y=215765
X1029 441 955 435 483 956 1 2 DFCND2BWP7T $T=387920 208160 0 0 $X=387630 $Y=207925
X1030 143 1 149 145 842 2 OAI21D2BWP7T $T=135360 208160 1 180 $X=130030 $Y=207925
X1031 146 1 159 157 808 2 OAI21D2BWP7T $T=142080 200320 1 180 $X=136750 $Y=200085
X1032 384 1 876 378 927 2 OAI21D2BWP7T $T=307280 216000 1 180 $X=301950 $Y=215765
X1033 442 423 1 438 944 2 IOA21D1BWP7T $T=361600 216000 1 180 $X=357950 $Y=215765
X1034 828 114 1 108 2 836 44 OAI22D1BWP7T $T=104560 216000 0 0 $X=104270 $Y=215765
X1035 790 845 1 130 2 854 839 OAI22D1BWP7T $T=135360 223840 1 180 $X=131150 $Y=223605
X1036 908 345 1 343 2 339 918 OAI22D1BWP7T $T=280960 223840 1 180 $X=276750 $Y=223605
X1037 934 345 1 343 2 413 935 OAI22D1BWP7T $T=335280 216000 0 0 $X=334990 $Y=215765
X1038 957 345 1 343 2 500 958 OAI22D1BWP7T $T=416480 223840 0 0 $X=416190 $Y=223605
X1039 220 862 220 197 223 1 2 225 AO221D1BWP7T $T=184640 216000 0 0 $X=184350 $Y=215765
X1040 365 369 356 921 357 1 2 374 AO221D1BWP7T $T=295520 216000 1 0 $X=295230 $Y=211790
X1041 392 396 397 398 400 1 2 403 AO221D1BWP7T $T=314000 208160 1 0 $X=313710 $Y=203950
X1042 536 538 540 967 456 1 2 547 AO221D1BWP7T $T=459040 223840 0 0 $X=458750 $Y=223605
X1043 537 458 965 964 456 1 2 546 AO221D1BWP7T $T=461280 223840 1 0 $X=460990 $Y=219630
X1044 214 311 208 907 2 1 906 DFCND0BWP7T $T=263600 200320 1 180 $X=250430 $Y=200085
X1045 214 910 208 915 2 1 326 DFCND0BWP7T $T=259120 231680 1 0 $X=258830 $Y=227470
X1046 214 913 208 321 2 1 270 DFCND0BWP7T $T=278160 200320 1 180 $X=264990 $Y=200085
X1047 441 950 435 968 2 1 467 DFCND0BWP7T $T=376720 216000 0 0 $X=376430 $Y=215765
X1048 441 954 435 969 2 1 480 DFCND0BWP7T $T=381200 208160 1 0 $X=380910 $Y=203950
X1049 324 306 322 320 316 314 2 912 1 OA222D0BWP7T $T=268640 208160 0 180 $X=262190 $Y=203950
X1050 916 306 234 915 316 321 2 911 1 OA222D0BWP7T $T=272000 216000 0 180 $X=265550 $Y=211790
X1051 327 306 234 325 316 323 2 909 1 OA222D0BWP7T $T=272560 223840 0 180 $X=266110 $Y=219630
X1052 306 917 1 234 915 316 318 2 910 OAI222D2BWP7T $T=273680 223840 1 180 $X=263310 $Y=223605
X1053 264 892 258 1 2 XOR2D2BWP7T $T=223280 216000 1 180 $X=216270 $Y=215765
X1054 178 228 237 239 2 1 IAO21D2BWP7T $T=194160 208160 0 0 $X=193870 $Y=207925
X1055 17 15 775 1 2 ND2D1P5BWP7T $T=27840 231680 0 180 $X=23630 $Y=227470
X1056 858 2 171 176 1 180 862 AOI211XD2BWP7T $T=142640 223840 0 0 $X=142350 $Y=223605
X1057 362 453 917 949 456 459 1 2 AO221D2BWP7T $T=375040 208160 0 0 $X=374750 $Y=207925
X1058 535 503 966 904 456 541 1 2 AO221D2BWP7T $T=457920 208160 1 0 $X=457630 $Y=203950
X1059 178 1 181 858 173 175 2 OAI22D2BWP7T $T=153280 223840 0 180 $X=146270 $Y=219630
X1060 178 1 181 855 173 175 2 OAI22D2BWP7T $T=156080 216000 0 180 $X=149070 $Y=211790
X1061 959 1 345 507 961 343 2 OAI22D2BWP7T $T=422640 223840 1 0 $X=422350 $Y=219630
X1062 179 2 169 855 1 172 NR3D3BWP7T $T=152160 208160 1 180 $X=140110 $Y=207925
X1063 860 263 896 860 2 263 1 IOA22D2BWP7T $T=227200 231680 0 180 $X=220750 $Y=227470
X1064 233 306 1 2 CKND8BWP7T $T=254080 216000 0 0 $X=253790 $Y=215765
X1065 187 2 178 1 244 NR2XD3BWP7T $T=189120 231680 1 0 $X=188830 $Y=227470
X1066 218 879 214 208 866 190 1 2 EDFCND2BWP7T $T=185200 223840 0 180 $X=166430 $Y=219630
X1067 150 2 158 168 861 860 1 NR4D4BWP7T $T=132560 208160 1 0 $X=132270 $Y=203950
X1068 829 1 823 2 833 OR2D0BWP7T $T=105680 216000 1 0 $X=105390 $Y=211790
X1069 70 1 67 54 794 2 793 IIND4D0BWP7T $T=67040 208160 0 180 $X=61710 $Y=203950
X1070 818 1 96 4 816 2 11 IIND4D0BWP7T $T=93920 208160 0 180 $X=88590 $Y=203950
X1071 93 90 803 67 2 85 1 IINR4D1BWP7T $T=91680 208160 1 180 $X=84110 $Y=207925
.ENDS
***************************************
.SUBCKT NR2D5BWP7T A2 VDD A1 VSS ZN
** N=6 EP=5 IP=0 FDC=20
M0 VSS A2 ZN VSS N L=1.8e-07 W=1e-06 $X=640 $Y=345 $D=0
M1 ZN A2 VSS VSS N L=1.8e-07 W=1e-06 $X=1420 $Y=345 $D=0
M2 VSS A2 ZN VSS N L=1.8e-07 W=1e-06 $X=2180 $Y=345 $D=0
M3 ZN A2 VSS VSS N L=1.8e-07 W=1e-06 $X=2920 $Y=345 $D=0
M4 VSS A2 ZN VSS N L=1.8e-07 W=1e-06 $X=3680 $Y=345 $D=0
M5 ZN A1 VSS VSS N L=1.8e-07 W=1e-06 $X=4440 $Y=345 $D=0
M6 VSS A1 ZN VSS N L=1.8e-07 W=1e-06 $X=5200 $Y=345 $D=0
M7 ZN A1 VSS VSS N L=1.8e-07 W=1e-06 $X=5940 $Y=345 $D=0
M8 VSS A1 ZN VSS N L=1.8e-07 W=1e-06 $X=6700 $Y=345 $D=0
M9 ZN A1 VSS VSS N L=1.8e-07 W=1e-06 $X=7480 $Y=345 $D=0
M10 6 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=640 $Y=2205 $D=16
M11 VDD A2 6 VDD P L=1.8e-07 W=1.37e-06 $X=1400 $Y=2205 $D=16
M12 6 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2160 $Y=2205 $D=16
M13 VDD A2 6 VDD P L=1.8e-07 W=1.37e-06 $X=2920 $Y=2205 $D=16
M14 6 A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3680 $Y=2205 $D=16
M15 ZN A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=4440 $Y=2205 $D=16
M16 6 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=5200 $Y=2205 $D=16
M17 ZN A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=5960 $Y=2205 $D=16
M18 6 A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=6720 $Y=2205 $D=16
M19 ZN A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=7480 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT INR2XD4BWP7T B1 ZN A1 VSS VDD
** N=7 EP=5 IP=0 FDC=32
M0 ZN B1 VSS VSS N L=1.8e-07 W=5.7e-07 $X=620 $Y=345 $D=0
M1 VSS B1 ZN VSS N L=1.8e-07 W=5.7e-07 $X=1340 $Y=345 $D=0
M2 ZN B1 VSS VSS N L=1.8e-07 W=5.7e-07 $X=2060 $Y=345 $D=0
M3 VSS B1 ZN VSS N L=1.8e-07 W=5.7e-07 $X=2780 $Y=345 $D=0
M4 ZN B1 VSS VSS N L=1.8e-07 W=5.7e-07 $X=3500 $Y=345 $D=0
M5 VSS B1 ZN VSS N L=1.8e-07 W=5.7e-07 $X=4220 $Y=345 $D=0
M6 ZN B1 VSS VSS N L=1.8e-07 W=5.7e-07 $X=4940 $Y=345 $D=0
M7 VSS 7 ZN VSS N L=1.8e-07 W=5.7e-07 $X=5660 $Y=345 $D=0
M8 ZN 7 VSS VSS N L=1.8e-07 W=5.7e-07 $X=6380 $Y=345 $D=0
M9 VSS 7 ZN VSS N L=1.8e-07 W=5.7e-07 $X=7100 $Y=345 $D=0
M10 ZN 7 VSS VSS N L=1.8e-07 W=5.7e-07 $X=7820 $Y=345 $D=0
M11 VSS 7 ZN VSS N L=1.8e-07 W=5.7e-07 $X=8540 $Y=345 $D=0
M12 ZN 7 VSS VSS N L=1.8e-07 W=5.7e-07 $X=9260 $Y=345 $D=0
M13 VSS 7 ZN VSS N L=1.8e-07 W=5.7e-07 $X=9980 $Y=345 $D=0
M14 7 A1 VSS VSS N L=1.8e-07 W=1e-06 $X=11360 $Y=345 $D=0
M15 VSS A1 7 VSS N L=1.8e-07 W=1e-06 $X=12080 $Y=345 $D=0
M16 6 B1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M17 VDD B1 6 VDD P L=1.8e-07 W=1.555e-06 $X=1340 $Y=2020 $D=16
M18 6 B1 VDD VDD P L=1.8e-07 W=1.555e-06 $X=2060 $Y=2020 $D=16
M19 VDD B1 6 VDD P L=1.8e-07 W=1.555e-06 $X=2780 $Y=2020 $D=16
M20 6 B1 VDD VDD P L=1.8e-07 W=1.555e-06 $X=3500 $Y=2020 $D=16
M21 VDD B1 6 VDD P L=1.8e-07 W=1.555e-06 $X=4220 $Y=2020 $D=16
M22 6 B1 VDD VDD P L=1.8e-07 W=1.555e-06 $X=4940 $Y=2020 $D=16
M23 ZN 7 6 VDD P L=1.8e-07 W=1.555e-06 $X=5660 $Y=2020 $D=16
M24 6 7 ZN VDD P L=1.8e-07 W=1.555e-06 $X=6380 $Y=2020 $D=16
M25 ZN 7 6 VDD P L=1.8e-07 W=1.555e-06 $X=7100 $Y=2020 $D=16
M26 6 7 ZN VDD P L=1.8e-07 W=1.555e-06 $X=7820 $Y=2020 $D=16
M27 ZN 7 6 VDD P L=1.8e-07 W=1.555e-06 $X=8540 $Y=2020 $D=16
M28 6 7 ZN VDD P L=1.8e-07 W=1.555e-06 $X=9260 $Y=2020 $D=16
M29 ZN 7 6 VDD P L=1.8e-07 W=1.37e-06 $X=9980 $Y=2205 $D=16
M30 7 A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=11360 $Y=2205 $D=16
M31 VDD A1 7 VDD P L=1.8e-07 W=1.37e-06 $X=12080 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT OR2D1BWP7T A1 VSS A2 VDD Z
** N=7 EP=5 IP=0 FDC=6
M0 6 A1 VSS VSS N L=1.8e-07 W=5e-07 $X=660 $Y=845 $D=0
M1 VSS A2 6 VSS N L=1.8e-07 W=5e-07 $X=1380 $Y=845 $D=0
M2 Z 6 VSS VSS N L=1.8e-07 W=1e-06 $X=2000 $Y=345 $D=0
M3 7 A1 6 VDD P L=1.8e-07 W=1.37e-06 $X=660 $Y=2205 $D=16
M4 VDD A2 7 VDD P L=1.8e-07 W=1.37e-06 $X=1200 $Y=2205 $D=16
M5 Z 6 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2000 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300 301
+ 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321
+ 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341
+ 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361
+ 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381
+ 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401
+ 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421
+ 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441
+ 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461
+ 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481
+ 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501
+ 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521
+ 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541
+ 542 543 544
** N=934 EP=543 IP=3729 FDC=4877
M0 926 214 1 1 N L=1.8e-07 W=5e-07 $X=197620 $Y=191535 $D=0
M1 841 194 926 1 N L=1.8e-07 W=5e-07 $X=198260 $Y=191535 $D=0
M2 927 841 1 1 N L=1.8e-07 W=1e-06 $X=207875 $Y=192825 $D=0
M3 928 834 927 1 N L=1.8e-07 W=1e-06 $X=208725 $Y=192825 $D=0
M4 929 842 928 1 N L=1.8e-07 W=1e-06 $X=209570 $Y=192825 $D=0
M5 848 257 929 1 N L=1.8e-07 W=1e-06 $X=210430 $Y=192825 $D=0
M6 930 257 848 1 N L=1.8e-07 W=1e-06 $X=211300 $Y=192825 $D=0
M7 931 842 930 1 N L=1.8e-07 W=1e-06 $X=211985 $Y=192825 $D=0
M8 932 834 931 1 N L=1.8e-07 W=1e-06 $X=212670 $Y=192825 $D=0
M9 1 841 932 1 N L=1.8e-07 W=1e-06 $X=213355 $Y=192825 $D=0
M10 261 848 1 1 N L=1.8e-07 W=1e-06 $X=214160 $Y=192825 $D=0
M11 1 848 261 1 N L=1.8e-07 W=1e-06 $X=214880 $Y=192825 $D=0
M12 261 848 1 1 N L=1.8e-07 W=1e-06 $X=215600 $Y=192825 $D=0
M13 1 848 261 1 N L=1.8e-07 W=1e-06 $X=216320 $Y=192825 $D=0
M14 933 327 907 1 N L=1.8e-07 W=1e-06 $X=361100 $Y=184985 $D=0
M15 1 410 933 1 N L=1.8e-07 W=1e-06 $X=361645 $Y=184985 $D=0
M16 934 326 1 1 N L=1.8e-07 W=1e-06 $X=362540 $Y=184985 $D=0
M17 907 414 934 1 N L=1.8e-07 W=1e-06 $X=363025 $Y=184985 $D=0
M18 417 907 1 1 N L=1.8e-07 W=1e-06 $X=364545 $Y=184985 $D=0
M19 1 907 417 1 N L=1.8e-07 W=1e-06 $X=365280 $Y=184985 $D=0
M20 841 214 2 2 P L=1.8e-07 W=6.85e-07 $X=197620 $Y=189165 $D=16
M21 2 194 841 2 P L=1.8e-07 W=6.85e-07 $X=198340 $Y=189165 $D=16
M22 848 841 2 2 P L=1.8e-07 W=1.37e-06 $X=207875 $Y=194685 $D=16
M23 2 834 848 2 P L=1.8e-07 W=1.37e-06 $X=208600 $Y=194685 $D=16
M24 848 842 2 2 P L=1.8e-07 W=1.305e-06 $X=209570 $Y=194750 $D=16
M25 2 257 848 2 P L=1.8e-07 W=1.305e-06 $X=210400 $Y=194750 $D=16
M26 848 257 2 2 P L=1.8e-07 W=1.305e-06 $X=211200 $Y=194750 $D=16
M27 2 842 848 2 P L=1.8e-07 W=1.305e-06 $X=211920 $Y=194750 $D=16
M28 848 834 2 2 P L=1.8e-07 W=1.37e-06 $X=212720 $Y=194685 $D=16
M29 2 841 848 2 P L=1.8e-07 W=1.37e-06 $X=213440 $Y=194685 $D=16
M30 261 848 2 2 P L=1.8e-07 W=1.37e-06 $X=214160 $Y=194685 $D=16
M31 2 848 261 2 P L=1.8e-07 W=1.37e-06 $X=214880 $Y=194685 $D=16
M32 261 848 2 2 P L=1.8e-07 W=1.37e-06 $X=215600 $Y=194685 $D=16
M33 2 848 261 2 P L=1.8e-07 W=1.37e-06 $X=216320 $Y=194685 $D=16
M34 2 327 906 2 P L=1.8e-07 W=1.37e-06 $X=361100 $Y=186845 $D=16
M35 906 410 2 2 P L=1.8e-07 W=1.37e-06 $X=361820 $Y=186845 $D=16
M36 907 326 906 2 P L=1.8e-07 W=1.37e-06 $X=362540 $Y=186845 $D=16
M37 906 414 907 2 P L=1.8e-07 W=1.37e-06 $X=363260 $Y=186845 $D=16
M38 417 907 2 2 P L=1.8e-07 W=1.37e-06 $X=364545 $Y=186845 $D=16
M39 2 907 417 2 P L=1.8e-07 W=1.37e-06 $X=365280 $Y=186845 $D=16
X102 1 500 ANTENNABWP7T $T=470800 200320 0 180 $X=469390 $Y=196110
X103 1 532 ANTENNABWP7T $T=470800 168960 0 0 $X=470510 $Y=168725
X104 1 534 ANTENNABWP7T $T=471920 176800 0 180 $X=470510 $Y=172590
X105 1 343 ANTENNABWP7T $T=470800 176800 0 0 $X=470510 $Y=176565
X106 1 535 ANTENNABWP7T $T=471920 184640 0 180 $X=470510 $Y=180430
X107 1 360 ANTENNABWP7T $T=470800 184640 0 0 $X=470510 $Y=184405
X108 1 480 ANTENNABWP7T $T=471920 192480 0 180 $X=470510 $Y=188270
X109 1 533 ANTENNABWP7T $T=470800 192480 0 0 $X=470510 $Y=192245
X110 1 527 ANTENNABWP7T $T=471920 200320 0 180 $X=470510 $Y=196110
X111 1 536 ANTENNABWP7T $T=471920 168960 0 0 $X=471630 $Y=168725
X112 1 537 ANTENNABWP7T $T=473040 176800 0 180 $X=471630 $Y=172590
X113 1 495 ANTENNABWP7T $T=471920 176800 0 0 $X=471630 $Y=176565
X114 1 488 ANTENNABWP7T $T=473040 184640 0 180 $X=471630 $Y=180430
X115 1 518 ANTENNABWP7T $T=471920 184640 0 0 $X=471630 $Y=184405
X116 1 538 ANTENNABWP7T $T=473040 192480 0 180 $X=471630 $Y=188270
X117 1 531 ANTENNABWP7T $T=471920 192480 0 0 $X=471630 $Y=192245
X118 1 539 ANTENNABWP7T $T=473040 200320 0 180 $X=471630 $Y=196110
X119 1 544 ANTENNABWP7T $T=473040 168960 0 0 $X=472750 $Y=168725
X120 1 330 ANTENNABWP7T $T=474160 176800 0 180 $X=472750 $Y=172590
X121 1 540 ANTENNABWP7T $T=473040 176800 0 0 $X=472750 $Y=176565
X122 1 542 ANTENNABWP7T $T=474160 184640 0 180 $X=472750 $Y=180430
X123 1 439 ANTENNABWP7T $T=473040 184640 0 0 $X=472750 $Y=184405
X124 1 474 ANTENNABWP7T $T=474160 192480 0 180 $X=472750 $Y=188270
X125 1 541 ANTENNABWP7T $T=473040 192480 0 0 $X=472750 $Y=192245
X126 1 543 ANTENNABWP7T $T=474160 200320 0 180 $X=472750 $Y=196110
X184 808 1 2 181 CKBD1BWP7T $T=146560 176800 1 180 $X=144030 $Y=176565
X185 823 1 2 253 CKBD1BWP7T $T=206480 184640 0 0 $X=206190 $Y=184405
X186 879 1 2 310 CKBD1BWP7T $T=266400 184640 1 0 $X=266110 $Y=180430
X187 330 1 2 329 CKBD1BWP7T $T=292160 176800 1 180 $X=289630 $Y=176565
X188 900 1 2 375 CKBD1BWP7T $T=325200 200320 0 180 $X=322670 $Y=196110
X189 908 1 2 415 CKBD1BWP7T $T=366640 192480 1 180 $X=364110 $Y=192245
X190 439 1 2 425 CKBD1BWP7T $T=389040 176800 1 180 $X=386510 $Y=176565
X191 913 1 2 463 CKBD1BWP7T $T=403600 200320 1 0 $X=403310 $Y=196110
X192 480 1 2 916 CKBD1BWP7T $T=423200 192480 0 0 $X=422910 $Y=192245
X193 488 1 2 431 CKBD1BWP7T $T=432720 184640 1 180 $X=430190 $Y=184405
X194 492 1 2 493 CKBD1BWP7T $T=430480 192480 0 0 $X=430190 $Y=192245
X195 500 1 2 492 CKBD1BWP7T $T=440000 192480 0 180 $X=437470 $Y=188270
X196 43 1 2 763 INVD0BWP7T $T=44080 200320 0 180 $X=42110 $Y=196110
X197 57 1 2 59 INVD0BWP7T $T=51360 168960 0 0 $X=51070 $Y=168725
X198 761 1 2 775 INVD0BWP7T $T=68720 184640 0 0 $X=68430 $Y=184405
X199 41 1 2 91 INVD0BWP7T $T=80480 168960 0 0 $X=80190 $Y=168725
X200 65 1 2 114 INVD0BWP7T $T=92800 192480 0 0 $X=92510 $Y=192245
X201 119 1 2 108 INVD0BWP7T $T=97840 168960 1 180 $X=95870 $Y=168725
X202 68 1 2 123 INVD0BWP7T $T=98960 168960 0 0 $X=98670 $Y=168725
X203 113 1 2 161 INVD0BWP7T $T=128640 200320 0 180 $X=126670 $Y=196110
X204 222 1 2 238 INVD0BWP7T $T=182960 176800 1 0 $X=182670 $Y=172590
X205 861 1 2 857 INVD0BWP7T $T=226080 176800 1 0 $X=225790 $Y=172590
X206 855 1 2 866 INVD0BWP7T $T=230000 192480 0 0 $X=229710 $Y=192245
X207 283 1 2 875 INVD0BWP7T $T=247920 184640 1 0 $X=247630 $Y=180430
X208 882 1 2 881 INVD0BWP7T $T=270880 192480 0 180 $X=268910 $Y=188270
X209 884 1 2 883 INVD0BWP7T $T=274240 176800 1 180 $X=272270 $Y=176565
X210 330 1 2 890 INVD0BWP7T $T=293840 176800 1 180 $X=291870 $Y=176565
X211 328 1 2 886 INVD0BWP7T $T=294960 192480 0 180 $X=292990 $Y=188270
X212 332 1 2 891 INVD0BWP7T $T=296080 200320 0 180 $X=294110 $Y=196110
X213 274 1 2 895 INVD0BWP7T $T=306720 192480 0 180 $X=304750 $Y=188270
X214 856 1 2 894 INVD0BWP7T $T=305600 176800 0 0 $X=305310 $Y=176565
X215 368 1 2 896 INVD0BWP7T $T=315120 176800 0 180 $X=313150 $Y=172590
X216 860 1 2 899 INVD0BWP7T $T=317920 168960 0 0 $X=317630 $Y=168725
X217 364 1 2 897 INVD0BWP7T $T=320160 200320 0 180 $X=318190 $Y=196110
X218 406 1 2 905 INVD0BWP7T $T=359360 168960 1 180 $X=357390 $Y=168725
X219 420 1 2 911 INVD0BWP7T $T=387920 184640 1 180 $X=385950 $Y=184405
X220 449 1 2 912 INVD0BWP7T $T=395200 168960 0 0 $X=394910 $Y=168725
X221 488 1 2 489 INVD0BWP7T $T=428240 168960 0 0 $X=427950 $Y=168725
X222 494 1 2 918 INVD0BWP7T $T=434400 184640 0 0 $X=434110 $Y=184405
X223 496 1 2 917 INVD0BWP7T $T=434960 200320 1 0 $X=434670 $Y=196110
X224 479 1 2 922 INVD0BWP7T $T=437760 176800 0 0 $X=437470 $Y=176565
X225 500 1 2 502 INVD0BWP7T $T=440000 192480 1 0 $X=439710 $Y=188270
X226 316 1 2 919 INVD0BWP7T $T=442800 184640 1 180 $X=440830 $Y=184405
X227 509 1 2 923 INVD0BWP7T $T=443920 192480 1 0 $X=443630 $Y=188270
X228 501 1 2 921 INVD0BWP7T $T=451200 192480 1 180 $X=449230 $Y=192245
X229 516 1 2 925 INVD0BWP7T $T=461280 192480 0 0 $X=460990 $Y=192245
X230 486 1 2 924 INVD0BWP7T $T=465760 192480 1 180 $X=463790 $Y=192245
X231 830 256 1 2 BUFFD1P5BWP7T $T=207040 176800 1 0 $X=206750 $Y=172590
X232 822 266 1 2 BUFFD1P5BWP7T $T=218800 168960 0 0 $X=218510 $Y=168725
X233 360 357 1 2 BUFFD1P5BWP7T $T=313440 192480 1 180 $X=310350 $Y=192245
X234 495 498 1 2 BUFFD1P5BWP7T $T=434400 176800 0 0 $X=434110 $Y=176565
X235 504 856 1 2 BUFFD1P5BWP7T $T=442800 192480 1 180 $X=439710 $Y=192245
X236 518 860 1 2 BUFFD1P5BWP7T $T=463520 184640 0 180 $X=460430 $Y=180430
X237 527 316 1 2 BUFFD1P5BWP7T $T=468560 184640 1 180 $X=465470 $Y=184405
X238 531 528 1 2 BUFFD1P5BWP7T $T=470800 192480 1 180 $X=467710 $Y=192245
X294 789 1 2 785 BUFFD1BWP7T $T=102880 168960 1 180 $X=100350 $Y=168725
X295 803 1 2 163 BUFFD1BWP7T $T=130880 176800 1 180 $X=128350 $Y=176565
X296 820 1 2 822 BUFFD1BWP7T $T=176240 168960 0 0 $X=175950 $Y=168725
X297 835 1 2 838 BUFFD1BWP7T $T=191360 176800 0 0 $X=191070 $Y=176565
X298 844 1 2 847 BUFFD1BWP7T $T=211520 176800 0 0 $X=211230 $Y=176565
X299 838 1 2 264 BUFFD1BWP7T $T=216560 168960 0 0 $X=216270 $Y=168725
X300 343 1 2 893 BUFFD1BWP7T $T=300560 176800 0 0 $X=300270 $Y=176565
X301 892 1 2 344 BUFFD1BWP7T $T=303920 192480 1 180 $X=301390 $Y=192245
X302 362 1 2 359 BUFFD1BWP7T $T=314000 168960 1 180 $X=311470 $Y=168725
X303 405 1 2 904 BUFFD1BWP7T $T=359360 200320 0 180 $X=356830 $Y=196110
X304 909 1 2 418 BUFFD1BWP7T $T=374480 184640 1 0 $X=374190 $Y=180430
X305 420 1 2 910 BUFFD1BWP7T $T=375040 184640 0 0 $X=374750 $Y=184405
X306 431 1 2 429 BUFFD1BWP7T $T=381760 200320 0 180 $X=379230 $Y=196110
X307 914 1 2 468 BUFFD1BWP7T $T=406960 184640 0 0 $X=406670 $Y=184405
X308 401 1 2 471 BUFFD1BWP7T $T=415920 192480 0 0 $X=415630 $Y=192245
X309 920 1 2 506 BUFFD1BWP7T $T=441120 184640 1 0 $X=440830 $Y=180430
X310 510 1 2 511 BUFFD1BWP7T $T=443920 200320 1 0 $X=443630 $Y=196110
X311 529 1 2 530 BUFFD1BWP7T $T=467440 200320 1 0 $X=467150 $Y=196110
X312 1 2 DCAP4BWP7T $T=55280 184640 1 0 $X=54990 $Y=180430
X313 1 2 DCAP4BWP7T $T=67040 176800 0 0 $X=66750 $Y=176565
X314 1 2 DCAP4BWP7T $T=135360 168960 0 0 $X=135070 $Y=168725
X315 1 2 DCAP4BWP7T $T=136480 176800 0 0 $X=136190 $Y=176565
X316 1 2 DCAP4BWP7T $T=143760 176800 1 0 $X=143470 $Y=172590
X317 1 2 DCAP4BWP7T $T=203120 168960 0 0 $X=202830 $Y=168725
X318 1 2 DCAP4BWP7T $T=226080 200320 1 0 $X=225790 $Y=196110
X319 1 2 DCAP4BWP7T $T=226640 184640 0 0 $X=226350 $Y=184405
X320 1 2 DCAP4BWP7T $T=227760 192480 0 0 $X=227470 $Y=192245
X321 1 2 DCAP4BWP7T $T=235600 192480 1 0 $X=235310 $Y=188270
X322 1 2 DCAP4BWP7T $T=241760 176800 0 0 $X=241470 $Y=176565
X323 1 2 DCAP4BWP7T $T=250720 176800 1 0 $X=250430 $Y=172590
X324 1 2 DCAP4BWP7T $T=283760 200320 1 0 $X=283470 $Y=196110
X325 1 2 DCAP4BWP7T $T=413120 176800 1 0 $X=412830 $Y=172590
X326 1 2 DCAP4BWP7T $T=422080 192480 1 0 $X=421790 $Y=188270
X327 1 2 DCAP4BWP7T $T=435520 192480 1 0 $X=435230 $Y=188270
X328 1 2 DCAP4BWP7T $T=451760 184640 0 0 $X=451470 $Y=184405
X329 1 2 DCAP4BWP7T $T=468560 184640 0 0 $X=468270 $Y=184405
X330 1 2 ICV_3 $T=31200 176800 0 0 $X=30910 $Y=176565
X331 1 2 ICV_3 $T=35120 184640 1 0 $X=34830 $Y=180430
X332 1 2 ICV_3 $T=35120 200320 1 0 $X=34830 $Y=196110
X333 1 2 ICV_3 $T=44640 176800 1 0 $X=44350 $Y=172590
X334 1 2 ICV_3 $T=53040 176800 0 0 $X=52750 $Y=176565
X335 1 2 ICV_3 $T=55280 192480 1 0 $X=54990 $Y=188270
X336 1 2 ICV_3 $T=65360 176800 1 0 $X=65070 $Y=172590
X337 1 2 ICV_3 $T=77120 192480 0 0 $X=76830 $Y=192245
X338 1 2 ICV_3 $T=88880 200320 1 0 $X=88590 $Y=196110
X339 1 2 ICV_3 $T=115200 192480 0 0 $X=114910 $Y=192245
X340 1 2 ICV_3 $T=119120 168960 0 0 $X=118830 $Y=168725
X341 1 2 ICV_3 $T=119120 184640 1 0 $X=118830 $Y=180430
X342 1 2 ICV_3 $T=119120 192480 1 0 $X=118830 $Y=188270
X343 1 2 ICV_3 $T=119120 200320 1 0 $X=118830 $Y=196110
X344 1 2 ICV_3 $T=145440 200320 1 0 $X=145150 $Y=196110
X345 1 2 ICV_3 $T=149920 168960 0 0 $X=149630 $Y=168725
X346 1 2 ICV_3 $T=157200 176800 1 0 $X=156910 $Y=172590
X347 1 2 ICV_3 $T=157200 184640 1 0 $X=156910 $Y=180430
X348 1 2 ICV_3 $T=157200 184640 0 0 $X=156910 $Y=184405
X349 1 2 ICV_3 $T=161120 168960 0 0 $X=160830 $Y=168725
X350 1 2 ICV_3 $T=161120 176800 1 0 $X=160830 $Y=172590
X351 1 2 ICV_3 $T=161120 176800 0 0 $X=160830 $Y=176565
X352 1 2 ICV_3 $T=161120 184640 0 0 $X=160830 $Y=184405
X353 1 2 ICV_3 $T=161120 192480 0 0 $X=160830 $Y=192245
X354 1 2 ICV_3 $T=178480 184640 0 0 $X=178190 $Y=184405
X355 1 2 ICV_3 $T=188560 176800 0 0 $X=188270 $Y=176565
X356 1 2 ICV_3 $T=199200 184640 0 0 $X=198910 $Y=184405
X357 1 2 ICV_3 $T=241200 168960 0 0 $X=240910 $Y=168725
X358 1 2 ICV_3 $T=241200 184640 0 0 $X=240910 $Y=184405
X359 1 2 ICV_3 $T=241200 192480 0 0 $X=240910 $Y=192245
X360 1 2 ICV_3 $T=283200 176800 0 0 $X=282910 $Y=176565
X361 1 2 ICV_3 $T=283200 184640 0 0 $X=282910 $Y=184405
X362 1 2 ICV_3 $T=283200 192480 1 0 $X=282910 $Y=188270
X363 1 2 ICV_3 $T=283200 192480 0 0 $X=282910 $Y=192245
X364 1 2 ICV_3 $T=287120 176800 0 0 $X=286830 $Y=176565
X365 1 2 ICV_3 $T=287120 184640 0 0 $X=286830 $Y=184405
X366 1 2 ICV_3 $T=291600 184640 1 0 $X=291310 $Y=180430
X367 1 2 ICV_3 $T=291600 200320 1 0 $X=291310 $Y=196110
X368 1 2 ICV_3 $T=301680 184640 1 0 $X=301390 $Y=180430
X369 1 2 ICV_3 $T=307280 176800 0 0 $X=306990 $Y=176565
X370 1 2 ICV_3 $T=310640 176800 1 0 $X=310350 $Y=172590
X371 1 2 ICV_3 $T=325200 176800 0 0 $X=324910 $Y=176565
X372 1 2 ICV_3 $T=325200 200320 1 0 $X=324910 $Y=196110
X373 1 2 ICV_3 $T=338080 168960 0 0 $X=337790 $Y=168725
X374 1 2 ICV_3 $T=345920 184640 1 0 $X=345630 $Y=180430
X375 1 2 ICV_3 $T=409200 168960 0 0 $X=408910 $Y=168725
X376 1 2 ICV_3 $T=409200 176800 1 0 $X=408910 $Y=172590
X377 1 2 ICV_3 $T=409200 184640 1 0 $X=408910 $Y=180430
X378 1 2 ICV_3 $T=409200 184640 0 0 $X=408910 $Y=184405
X379 1 2 ICV_3 $T=413120 192480 0 0 $X=412830 $Y=192245
X380 1 2 ICV_3 $T=437200 192480 0 0 $X=436910 $Y=192245
X381 1 2 ICV_3 $T=451200 192480 1 0 $X=450910 $Y=188270
X382 1 2 ICV_3 $T=451200 192480 0 0 $X=450910 $Y=192245
X383 1 2 ICV_3 $T=459600 168960 0 0 $X=459310 $Y=168725
X384 1 2 ICV_3 $T=459600 176800 1 0 $X=459310 $Y=172590
X385 1 2 ICV_3 $T=468000 184640 1 0 $X=467710 $Y=180430
X386 1 2 DCAP8BWP7T $T=29520 168960 0 0 $X=29230 $Y=168725
X387 1 2 DCAP8BWP7T $T=35120 176800 1 0 $X=34830 $Y=172590
X388 1 2 DCAP8BWP7T $T=35120 192480 1 0 $X=34830 $Y=188270
X389 1 2 DCAP8BWP7T $T=35120 192480 0 0 $X=34830 $Y=192245
X390 1 2 DCAP8BWP7T $T=40720 168960 0 0 $X=40430 $Y=168725
X391 1 2 DCAP8BWP7T $T=45200 192480 0 0 $X=44910 $Y=192245
X392 1 2 DCAP8BWP7T $T=59200 192480 0 0 $X=58910 $Y=192245
X393 1 2 DCAP8BWP7T $T=77120 176800 1 0 $X=76830 $Y=172590
X394 1 2 DCAP8BWP7T $T=82160 168960 0 0 $X=81870 $Y=168725
X395 1 2 DCAP8BWP7T $T=94480 192480 0 0 $X=94190 $Y=192245
X396 1 2 DCAP8BWP7T $T=107360 192480 0 0 $X=107070 $Y=192245
X397 1 2 DCAP8BWP7T $T=124160 168960 0 0 $X=123870 $Y=168725
X398 1 2 DCAP8BWP7T $T=132000 184640 0 0 $X=131710 $Y=184405
X399 1 2 DCAP8BWP7T $T=135920 200320 1 0 $X=135630 $Y=196110
X400 1 2 DCAP8BWP7T $T=140960 184640 1 0 $X=140670 $Y=180430
X401 1 2 DCAP8BWP7T $T=141520 168960 0 0 $X=141230 $Y=168725
X402 1 2 DCAP8BWP7T $T=152720 176800 1 0 $X=152430 $Y=172590
X403 1 2 DCAP8BWP7T $T=154400 192480 1 0 $X=154110 $Y=188270
X404 1 2 DCAP8BWP7T $T=154960 192480 0 0 $X=154670 $Y=192245
X405 1 2 DCAP8BWP7T $T=209840 176800 1 0 $X=209550 $Y=172590
X406 1 2 DCAP8BWP7T $T=217120 192480 0 0 $X=216830 $Y=192245
X407 1 2 DCAP8BWP7T $T=238400 200320 1 0 $X=238110 $Y=196110
X408 1 2 DCAP8BWP7T $T=239520 192480 1 0 $X=239230 $Y=188270
X409 1 2 DCAP8BWP7T $T=254640 176800 1 0 $X=254350 $Y=172590
X410 1 2 DCAP8BWP7T $T=259120 184640 0 0 $X=258830 $Y=184405
X411 1 2 DCAP8BWP7T $T=264160 192480 0 0 $X=263870 $Y=192245
X412 1 2 DCAP8BWP7T $T=266400 176800 1 0 $X=266110 $Y=172590
X413 1 2 DCAP8BWP7T $T=270880 192480 1 0 $X=270590 $Y=188270
X414 1 2 DCAP8BWP7T $T=278720 192480 1 0 $X=278430 $Y=188270
X415 1 2 DCAP8BWP7T $T=297200 184640 1 0 $X=296910 $Y=180430
X416 1 2 DCAP8BWP7T $T=297760 168960 0 0 $X=297470 $Y=168725
X417 1 2 DCAP8BWP7T $T=303920 192480 0 0 $X=303630 $Y=192245
X418 1 2 DCAP8BWP7T $T=306160 176800 1 0 $X=305870 $Y=172590
X419 1 2 DCAP8BWP7T $T=320720 176800 0 0 $X=320430 $Y=176565
X420 1 2 DCAP8BWP7T $T=322400 192480 0 0 $X=322110 $Y=192245
X421 1 2 DCAP8BWP7T $T=339760 200320 1 0 $X=339470 $Y=196110
X422 1 2 DCAP8BWP7T $T=341440 184640 1 0 $X=341150 $Y=180430
X423 1 2 DCAP8BWP7T $T=349840 200320 1 0 $X=349550 $Y=196110
X424 1 2 DCAP8BWP7T $T=352080 176800 0 0 $X=351790 $Y=176565
X425 1 2 DCAP8BWP7T $T=363840 168960 0 0 $X=363550 $Y=168725
X426 1 2 DCAP8BWP7T $T=363840 184640 1 0 $X=363550 $Y=180430
X427 1 2 DCAP8BWP7T $T=364960 176800 0 0 $X=364670 $Y=176565
X428 1 2 DCAP8BWP7T $T=381200 176800 0 0 $X=380910 $Y=176565
X429 1 2 DCAP8BWP7T $T=396880 168960 0 0 $X=396590 $Y=168725
X430 1 2 DCAP8BWP7T $T=401920 184640 0 0 $X=401630 $Y=184405
X431 1 2 DCAP8BWP7T $T=404720 184640 1 0 $X=404430 $Y=180430
X432 1 2 DCAP8BWP7T $T=405840 192480 1 0 $X=405550 $Y=188270
X433 1 2 DCAP8BWP7T $T=405840 200320 1 0 $X=405550 $Y=196110
X434 1 2 DCAP8BWP7T $T=422080 168960 0 0 $X=421790 $Y=168725
X435 1 2 DCAP8BWP7T $T=424880 184640 0 0 $X=424590 $Y=184405
X436 1 2 DCAP8BWP7T $T=463520 184640 1 0 $X=463230 $Y=180430
X437 2 1 DCAPBWP7T $T=21120 184640 0 0 $X=20830 $Y=184405
X438 2 1 DCAPBWP7T $T=25600 168960 0 0 $X=25310 $Y=168725
X439 2 1 DCAPBWP7T $T=32320 184640 0 0 $X=32030 $Y=184405
X440 2 1 DCAPBWP7T $T=41840 176800 0 0 $X=41550 $Y=176565
X441 2 1 DCAPBWP7T $T=45200 184640 1 0 $X=44910 $Y=180430
X442 2 1 DCAPBWP7T $T=84400 192480 0 0 $X=84110 $Y=192245
X443 2 1 DCAPBWP7T $T=125840 192480 0 0 $X=125550 $Y=192245
X444 2 1 DCAPBWP7T $T=140960 192480 1 0 $X=140670 $Y=188270
X445 2 1 DCAPBWP7T $T=167840 184640 0 0 $X=167550 $Y=184405
X446 2 1 DCAPBWP7T $T=174560 192480 1 0 $X=174270 $Y=188270
X447 2 1 DCAPBWP7T $T=192480 168960 0 0 $X=192190 $Y=168725
X448 2 1 DCAPBWP7T $T=209840 176800 0 0 $X=209550 $Y=176565
X449 2 1 DCAPBWP7T $T=242320 176800 1 0 $X=242030 $Y=172590
X450 2 1 DCAPBWP7T $T=251840 168960 0 0 $X=251550 $Y=168725
X451 2 1 DCAPBWP7T $T=276480 168960 0 0 $X=276190 $Y=168725
X452 2 1 DCAPBWP7T $T=284320 176800 1 0 $X=284030 $Y=172590
X453 2 1 DCAPBWP7T $T=303360 192480 1 0 $X=303070 $Y=188270
X454 2 1 DCAPBWP7T $T=326320 168960 0 0 $X=326030 $Y=168725
X455 2 1 DCAPBWP7T $T=335840 184640 0 0 $X=335550 $Y=184405
X456 2 1 DCAPBWP7T $T=335840 192480 0 0 $X=335550 $Y=192245
X457 2 1 DCAPBWP7T $T=338080 176800 0 0 $X=337790 $Y=176565
X458 2 1 DCAPBWP7T $T=356560 176800 0 0 $X=356270 $Y=176565
X459 2 1 DCAPBWP7T $T=368320 168960 0 0 $X=368030 $Y=168725
X460 2 1 DCAPBWP7T $T=368320 184640 1 0 $X=368030 $Y=180430
X461 2 1 DCAPBWP7T $T=368320 200320 1 0 $X=368030 $Y=196110
X462 2 1 DCAPBWP7T $T=399120 176800 1 0 $X=398830 $Y=172590
X463 2 1 DCAPBWP7T $T=410320 192480 1 0 $X=410030 $Y=188270
X464 2 1 DCAPBWP7T $T=410320 200320 1 0 $X=410030 $Y=196110
X465 2 1 DCAPBWP7T $T=426560 168960 0 0 $X=426270 $Y=168725
X466 2 1 DCAPBWP7T $T=432720 184640 0 0 $X=432430 $Y=184405
X467 2 1 DCAPBWP7T $T=433280 200320 1 0 $X=432990 $Y=196110
X468 2 1 DCAPBWP7T $T=443920 176800 0 0 $X=443630 $Y=176565
X469 2 1 DCAPBWP7T $T=452320 176800 0 0 $X=452030 $Y=176565
X470 2 1 DCAPBWP7T $T=452320 184640 1 0 $X=452030 $Y=180430
X471 274 381 383 326 368 327 1 2 903 AO222D0BWP7T $T=333600 192480 1 0 $X=333310 $Y=188270
X472 910 381 433 326 412 327 1 2 440 AO222D0BWP7T $T=382320 184640 1 0 $X=382030 $Y=180430
X473 486 381 483 326 479 327 1 2 476 AO222D0BWP7T $T=427680 176800 1 180 $X=421230 $Y=176565
X474 497 1 494 316 918 2 920 919 OAI221D1BWP7T $T=436080 184640 1 0 $X=435790 $Y=180430
X475 390 381 326 856 385 327 1 2 382 AO222D1BWP7T $T=341440 184640 0 180 $X=334430 $Y=180430
X476 462 381 326 455 453 327 1 2 450 AO222D1BWP7T $T=404720 184640 0 180 $X=397710 $Y=180430
X477 491 381 326 446 484 327 1 2 481 AO222D1BWP7T $T=431040 192480 0 180 $X=424030 $Y=188270
X478 490 381 326 487 485 327 1 2 482 AO222D1BWP7T $T=431600 176800 0 180 $X=424590 $Y=172590
X479 1 2 ICV_4 $T=21120 176800 0 0 $X=20830 $Y=176565
X480 1 2 ICV_4 $T=30080 184640 1 0 $X=29790 $Y=180430
X481 1 2 ICV_4 $T=114080 168960 0 0 $X=113790 $Y=168725
X482 1 2 ICV_4 $T=114080 192480 1 0 $X=113790 $Y=188270
X483 1 2 ICV_4 $T=203120 192480 0 0 $X=202830 $Y=192245
X484 1 2 ICV_4 $T=221600 168960 0 0 $X=221310 $Y=168725
X485 1 2 ICV_4 $T=222160 176800 1 0 $X=221870 $Y=172590
X486 1 2 ICV_4 $T=262480 184640 1 0 $X=262190 $Y=180430
X487 1 2 ICV_4 $T=274240 176800 0 0 $X=273950 $Y=176565
X488 1 2 ICV_4 $T=282080 184640 1 0 $X=281790 $Y=180430
X489 1 2 ICV_4 $T=287120 168960 0 0 $X=286830 $Y=168725
X490 1 2 ICV_4 $T=314000 168960 0 0 $X=313710 $Y=168725
X491 1 2 ICV_4 $T=324080 192480 1 0 $X=323790 $Y=188270
X492 1 2 ICV_4 $T=366080 184640 0 0 $X=365790 $Y=184405
X493 1 2 ICV_4 $T=371120 168960 0 0 $X=370830 $Y=168725
X494 1 2 ICV_4 $T=371120 184640 0 0 $X=370830 $Y=184405
X495 1 2 ICV_4 $T=455120 200320 1 0 $X=454830 $Y=196110
X496 400 903 393 2 1 342 DFCNQD1BWP7T $T=352080 176800 1 180 $X=339470 $Y=176565
X695 1 2 ICV_9 $T=20000 168960 0 0 $X=19710 $Y=168725
X696 1 2 ICV_9 $T=34000 176800 0 0 $X=33710 $Y=176565
X697 1 2 ICV_9 $T=34000 184640 0 0 $X=33710 $Y=184405
X698 1 2 ICV_9 $T=160000 184640 1 0 $X=159710 $Y=180430
X699 1 2 ICV_9 $T=202000 184640 1 0 $X=201710 $Y=180430
X700 1 2 ICV_9 $T=244000 176800 0 0 $X=243710 $Y=176565
X701 1 2 ICV_9 $T=244000 192480 1 0 $X=243710 $Y=188270
X702 1 2 ICV_9 $T=244000 192480 0 0 $X=243710 $Y=192245
X703 1 2 ICV_9 $T=286000 176800 1 0 $X=285710 $Y=172590
X704 1 2 ICV_9 $T=286000 184640 1 0 $X=285710 $Y=180430
X705 1 2 ICV_9 $T=286000 192480 1 0 $X=285710 $Y=188270
X706 1 2 ICV_9 $T=286000 192480 0 0 $X=285710 $Y=192245
X707 1 2 ICV_9 $T=286000 200320 1 0 $X=285710 $Y=196110
X708 1 2 ICV_9 $T=328000 184640 1 0 $X=327710 $Y=180430
X709 1 2 ICV_9 $T=328000 192480 1 0 $X=327710 $Y=188270
X710 1 2 ICV_9 $T=370000 192480 0 0 $X=369710 $Y=192245
X711 1 2 ICV_9 $T=370000 200320 1 0 $X=369710 $Y=196110
X712 1 2 ICV_9 $T=454000 168960 0 0 $X=453710 $Y=168725
X713 1 2 ICV_9 $T=454000 176800 1 0 $X=453710 $Y=172590
X714 1 2 ICV_9 $T=454000 184640 1 0 $X=453710 $Y=180430
X715 1 2 ICV_9 $T=454000 192480 1 0 $X=453710 $Y=188270
X716 1 2 ICV_9 $T=454000 192480 0 0 $X=453710 $Y=192245
X737 1 2 ICV_13 $T=30640 200320 1 0 $X=30350 $Y=196110
X738 1 2 ICV_13 $T=35120 168960 0 0 $X=34830 $Y=168725
X739 1 2 ICV_13 $T=72640 168960 0 0 $X=72350 $Y=168725
X740 1 2 ICV_13 $T=114640 184640 1 0 $X=114350 $Y=180430
X741 1 2 ICV_13 $T=130880 176800 1 0 $X=130590 $Y=172590
X742 1 2 ICV_13 $T=140960 176800 0 0 $X=140670 $Y=176565
X743 1 2 ICV_13 $T=161120 192480 1 0 $X=160830 $Y=188270
X744 1 2 ICV_13 $T=175120 184640 1 0 $X=174830 $Y=180430
X745 1 2 ICV_13 $T=182400 192480 1 0 $X=182110 $Y=188270
X746 1 2 ICV_13 $T=203120 184640 0 0 $X=202830 $Y=184405
X747 1 2 ICV_13 $T=245120 176800 1 0 $X=244830 $Y=172590
X748 1 2 ICV_13 $T=311200 192480 1 0 $X=310910 $Y=188270
X749 1 2 ICV_13 $T=324640 184640 1 0 $X=324350 $Y=180430
X750 1 2 ICV_13 $T=361040 192480 0 0 $X=360750 $Y=192245
X751 1 2 ICV_13 $T=366640 192480 0 0 $X=366350 $Y=192245
X752 1 2 ICV_13 $T=371120 184640 1 0 $X=370830 $Y=180430
X753 1 2 ICV_13 $T=400240 192480 0 0 $X=399950 $Y=192245
X754 1 2 ICV_13 $T=408640 192480 0 0 $X=408350 $Y=192245
X755 1 2 ICV_13 $T=432720 184640 1 0 $X=432430 $Y=180430
X756 372 373 2 373 898 372 1 MAOI22D1BWP7T $T=324080 192480 0 180 $X=319310 $Y=188270
X757 395 399 2 399 901 395 1 MAOI22D1BWP7T $T=353760 184640 1 180 $X=348990 $Y=184405
X758 12 1 2 6 INVD1BWP7T $T=23920 200320 0 180 $X=21950 $Y=196110
X759 757 1 2 20 INVD1BWP7T $T=27280 192480 1 180 $X=25310 $Y=192245
X760 18 1 2 759 INVD1BWP7T $T=27280 192480 1 0 $X=26990 $Y=188270
X761 58 1 2 3 INVD1BWP7T $T=53040 176800 1 180 $X=51070 $Y=176565
X762 788 1 2 16 INVD1BWP7T $T=99520 192480 0 0 $X=99230 $Y=192245
X763 157 1 2 175 INVD1BWP7T $T=137600 184640 0 0 $X=137310 $Y=184405
X764 847 1 2 876 INVD1BWP7T $T=252960 176800 1 0 $X=252670 $Y=172590
X765 322 1 2 320 INVD1BWP7T $T=278720 192480 0 180 $X=276750 $Y=188270
X766 331 1 2 334 INVD1BWP7T $T=292160 176800 1 0 $X=291870 $Y=172590
X767 339 1 2 335 INVD1BWP7T $T=296640 192480 0 180 $X=294670 $Y=188270
X768 338 1 2 319 INVD1BWP7T $T=296080 168960 0 0 $X=295790 $Y=168725
X769 387 1 2 388 INVD1BWP7T $T=339760 200320 0 180 $X=337790 $Y=196110
X770 408 1 2 411 INVD1BWP7T $T=360480 192480 1 0 $X=360190 $Y=188270
X771 421 1 2 422 INVD1BWP7T $T=378400 200320 0 180 $X=376430 $Y=196110
X772 451 1 2 452 INVD1BWP7T $T=398560 192480 0 0 $X=398270 $Y=192245
X773 471 1 2 469 INVD1BWP7T $T=418720 176800 0 180 $X=416750 $Y=172590
X774 1 2 DCAP16BWP7T $T=208160 192480 1 0 $X=207870 $Y=188270
X775 1 2 DCAP16BWP7T $T=217120 200320 1 0 $X=216830 $Y=196110
X776 1 2 DCAP16BWP7T $T=233360 176800 1 0 $X=233070 $Y=172590
X777 1 2 DCAP16BWP7T $T=274800 200320 1 0 $X=274510 $Y=196110
X778 1 2 DCAP16BWP7T $T=311760 176800 0 0 $X=311470 $Y=176565
X779 1 2 DCAP16BWP7T $T=329120 168960 0 0 $X=328830 $Y=168725
X780 1 2 DCAP16BWP7T $T=329120 176800 0 0 $X=328830 $Y=176565
X781 1 2 DCAP16BWP7T $T=329120 200320 1 0 $X=328830 $Y=196110
X782 1 2 DCAP16BWP7T $T=347600 168960 0 0 $X=347310 $Y=168725
X783 1 2 DCAP16BWP7T $T=359360 200320 1 0 $X=359070 $Y=196110
X784 1 2 DCAP16BWP7T $T=381200 192480 1 0 $X=380910 $Y=188270
X785 1 2 DCAP16BWP7T $T=381760 200320 1 0 $X=381470 $Y=196110
X786 1 2 DCAP16BWP7T $T=388480 184640 1 0 $X=388190 $Y=180430
X787 1 2 DCAP16BWP7T $T=390160 176800 1 0 $X=389870 $Y=172590
X788 1 2 DCAP16BWP7T $T=413120 192480 1 0 $X=412830 $Y=188270
X789 1 2 DCAP16BWP7T $T=423760 184640 1 0 $X=423470 $Y=180430
X790 1 2 DCAP16BWP7T $T=431600 176800 1 0 $X=431310 $Y=172590
X791 1 2 DCAP16BWP7T $T=442800 184640 0 0 $X=442510 $Y=184405
X792 1 2 DCAP16BWP7T $T=455120 184640 0 0 $X=454830 $Y=184405
X793 782 1 2 155 CKND1BWP7T $T=121920 200320 1 0 $X=121630 $Y=196110
X794 228 1 2 229 CKND1BWP7T $T=176800 192480 0 0 $X=176510 $Y=192245
X795 354 1 2 348 CKND1BWP7T $T=307840 200320 0 180 $X=305870 $Y=196110
X796 377 1 2 372 CKND1BWP7T $T=321840 168960 1 180 $X=319870 $Y=168725
X797 389 1 2 391 CKND1BWP7T $T=349840 200320 0 180 $X=347870 $Y=196110
X798 423 1 2 416 CKND1BWP7T $T=366640 176800 0 180 $X=364670 $Y=172590
X799 301 258 1 2 INVD4BWP7T $T=255760 200320 0 180 $X=251550 $Y=196110
X800 183 805 2 797 1 172 179 AOI22D1BWP7T $T=145440 200320 0 180 $X=141230 $Y=196110
X801 221 206 2 200 1 195 823 AOI22D1BWP7T $T=174560 184640 0 0 $X=174270 $Y=184405
X802 194 209 2 228 1 182 828 AOI22D1BWP7T $T=186880 200320 0 180 $X=182670 $Y=196110
X803 291 850 2 874 1 871 855 AOI22D1BWP7T $T=241200 192480 1 180 $X=236990 $Y=192245
X804 878 876 2 297 1 847 861 AOI22D1BWP7T $T=256320 176800 1 180 $X=252110 $Y=176565
X805 327 270 2 326 1 860 324 AOI22D1BWP7T $T=283200 192480 1 180 $X=278990 $Y=192245
X806 327 374 2 326 1 376 900 AOI22D1BWP7T $T=320720 184640 1 0 $X=320430 $Y=180430
X807 327 384 2 326 1 380 379 AOI22D1BWP7T $T=336400 176800 0 180 $X=332190 $Y=172590
X808 327 454 2 326 1 459 915 AOI22D1BWP7T $T=400800 176800 1 0 $X=400510 $Y=172590
X809 327 477 2 326 1 474 908 AOI22D1BWP7T $T=423760 184640 0 180 $X=419550 $Y=180430
X810 217 235 2 222 833 1 OAI21D1BWP7T $T=188000 176800 0 180 $X=184350 $Y=172590
X811 316 875 2 888 873 1 OAI21D1BWP7T $T=274240 184640 1 0 $X=273950 $Y=180430
X812 849 269 1 2 BUFFD8BWP7T $T=219360 176800 0 0 $X=219070 $Y=176565
X813 205 2 195 194 1 NR2D4BWP7T $T=157200 176800 1 180 $X=150190 $Y=176565
X814 849 265 1 2 BUFFD6BWP7T $T=215440 176800 1 0 $X=215150 $Y=172590
X815 470 428 1 2 BUFFD6BWP7T $T=418160 184640 0 0 $X=417870 $Y=184405
X816 33 23 2 1 INVD2BWP7T $T=38480 168960 0 0 $X=38190 $Y=168725
X817 171 758 2 1 INVD2BWP7T $T=138720 176800 0 0 $X=138430 $Y=176565
X818 204 209 2 1 INVD2BWP7T $T=163920 176800 0 0 $X=163630 $Y=176565
X819 398 397 2 1 INVD2BWP7T $T=350960 184640 0 180 $X=348430 $Y=180430
X820 261 403 2 1 INVD2BWP7T $T=381200 192480 0 180 $X=378670 $Y=188270
X821 446 442 2 1 INVD2BWP7T $T=392400 192480 1 180 $X=389870 $Y=192245
X822 467 466 2 1 INVD2BWP7T $T=409200 168960 1 180 $X=406670 $Y=168725
X823 503 508 2 1 INVD2BWP7T $T=447840 176800 1 180 $X=445310 $Y=176565
X824 515 517 2 1 INVD2BWP7T $T=462400 192480 0 180 $X=459870 $Y=188270
X825 852 856 1 2 859 CKXOR2D1BWP7T $T=221600 184640 1 0 $X=221310 $Y=180430
X826 877 876 1 2 298 CKXOR2D1BWP7T $T=259120 184640 1 180 $X=253790 $Y=184405
X827 847 885 1 2 889 CKXOR2D1BWP7T $T=278160 176800 0 0 $X=277870 $Y=176565
X828 889 330 1 2 887 CKXOR2D1BWP7T $T=291040 168960 0 0 $X=290750 $Y=168725
X829 270 854 152 1 2 CKXOR2D2BWP7T $T=227760 192480 1 180 $X=221310 $Y=192245
X830 904 401 396 1 2 CKXOR2D2BWP7T $T=355440 192480 0 180 $X=348990 $Y=188270
X831 2 1 DCAP32BWP7T $T=310080 184640 0 0 $X=309790 $Y=184405
X832 2 1 DCAP32BWP7T $T=343120 192480 0 0 $X=342830 $Y=192245
X833 160 802 162 71 1 2 OAI21D0BWP7T $T=130320 192480 0 180 $X=127230 $Y=188270
X834 207 808 205 212 1 2 OAI21D0BWP7T $T=163920 176800 1 0 $X=163630 $Y=172590
X835 193 813 209 202 1 2 OAI21D0BWP7T $T=167840 200320 1 0 $X=167550 $Y=196110
X836 221 218 217 816 1 2 OAI21D0BWP7T $T=171760 176800 1 180 $X=168670 $Y=176565
X837 243 837 193 182 1 2 OAI21D0BWP7T $T=193040 200320 0 180 $X=189950 $Y=196110
X838 857 868 860 858 1 2 OAI21D0BWP7T $T=228320 168960 0 0 $X=228030 $Y=168725
X839 865 863 274 280 1 2 OAI21D0BWP7T $T=231680 184640 0 0 $X=231390 $Y=184405
X840 866 872 284 276 1 2 OAI21D0BWP7T $T=235600 200320 1 0 $X=235310 $Y=196110
X841 434 436 437 276 1 2 OAI21D0BWP7T $T=385680 168960 0 0 $X=385390 $Y=168725
X842 272 851 1 2 852 XNR2D1BWP7T $T=230000 192480 0 180 $X=224670 $Y=188270
X843 120 122 2 1 CKND2BWP7T $T=97840 192480 1 0 $X=97550 $Y=188270
X844 186 806 2 1 CKND2BWP7T $T=148800 176800 1 180 $X=146270 $Y=176565
X845 200 190 2 1 CKND2BWP7T $T=154960 168960 1 180 $X=152430 $Y=168725
X846 201 243 2 1 CKND2BWP7T $T=195280 200320 0 180 $X=192750 $Y=196110
X847 207 831 2 1 CKND2BWP7T $T=196960 176800 1 0 $X=196670 $Y=172590
X848 270 323 2 1 CKND2BWP7T $T=277040 192480 0 0 $X=276750 $Y=192245
X849 472 475 2 1 CKND2BWP7T $T=419840 168960 0 0 $X=419550 $Y=168725
X850 210 1 2 816 CKND0BWP7T $T=165600 184640 1 0 $X=165310 $Y=180430
X851 850 1 2 871 CKND0BWP7T $T=239520 192480 0 180 $X=237550 $Y=188270
X852 356 1 2 358 CKND0BWP7T $T=310080 176800 0 0 $X=309790 $Y=176565
X853 412 1 2 413 CKND0BWP7T $T=362160 168960 0 0 $X=361870 $Y=168725
X854 831 2 205 826 814 180 1 AOI22D2BWP7T $T=188000 184640 1 180 $X=180990 $Y=184405
X855 227 2 833 842 831 205 1 AOI22D2BWP7T $T=189120 176800 1 0 $X=188830 $Y=172590
X856 288 2 850 865 871 286 1 AOI22D2BWP7T $T=241200 184640 1 180 $X=234190 $Y=184405
X857 299 2 876 281 847 302 1 AOI22D2BWP7T $T=253520 168960 0 0 $X=253230 $Y=168725
X858 327 2 353 349 352 326 1 AOI22D2BWP7T $T=311200 184640 0 180 $X=304190 $Y=180430
X859 327 2 369 363 359 326 1 AOI22D2BWP7T $T=320720 184640 0 180 $X=313710 $Y=180430
X860 327 2 409 902 407 326 1 AOI22D2BWP7T $T=364960 176800 1 180 $X=357950 $Y=176565
X861 327 2 438 432 435 326 1 AOI22D2BWP7T $T=390160 176800 0 180 $X=383150 $Y=172590
X862 327 2 478 473 916 326 1 AOI22D2BWP7T $T=426560 200320 0 180 $X=419550 $Y=196110
X863 233 230 180 200 199 2 1 AOI22D0BWP7T $T=176800 192480 1 180 $X=173150 $Y=192245
X864 342 892 290 327 326 2 1 AOI22D0BWP7T $T=298320 192480 0 0 $X=298030 $Y=192245
X865 347 345 893 327 326 2 1 AOI22D0BWP7T $T=303920 200320 0 180 $X=300270 $Y=196110
X866 199 1 2 810 CKBD0BWP7T $T=154960 192480 1 180 $X=152430 $Y=192245
X867 141 140 138 135 2 1 118 AO211D1BWP7T $T=110720 192480 0 180 $X=105950 $Y=188270
X868 22 2 13 16 1 NR2D1BWP7T $T=26160 200320 0 180 $X=23630 $Y=196110
X869 759 2 762 763 1 NR2D1BWP7T $T=28960 192480 1 0 $X=28670 $Y=188270
X870 779 2 89 88 1 NR2D1BWP7T $T=82160 192480 1 180 $X=79630 $Y=192245
X871 783 2 116 113 1 NR2D1BWP7T $T=91680 200320 1 0 $X=91390 $Y=196110
X872 95 2 126 127 1 NR2D1BWP7T $T=100640 176800 0 0 $X=100350 $Y=176565
X873 123 2 130 83 1 NR2D1BWP7T $T=103440 176800 1 0 $X=103150 $Y=172590
X874 109 2 141 152 1 NR2D1BWP7T $T=124160 168960 1 180 $X=121630 $Y=168725
X875 159 2 801 156 1 NR2D1BWP7T $T=126400 176800 0 0 $X=126110 $Y=176565
X876 204 2 811 182 1 NR2D1BWP7T $T=157200 184640 0 180 $X=154670 $Y=180430
X877 816 2 817 216 1 NR2D1BWP7T $T=166160 176800 0 0 $X=165870 $Y=176565
X878 235 2 814 206 1 NR2D1BWP7T $T=192480 184640 1 180 $X=189950 $Y=184405
X879 281 2 289 290 1 NR2D1BWP7T $T=238960 168960 0 0 $X=238670 $Y=168725
X880 847 2 870 293 1 NR2D1BWP7T $T=248480 176800 1 0 $X=248190 $Y=172590
X881 816 213 216 817 1 2 AOI21D0BWP7T $T=166720 176800 1 0 $X=166430 $Y=172590
X882 184 819 223 187 1 2 AOI21D0BWP7T $T=171200 168960 0 0 $X=170910 $Y=168725
X883 234 236 197 229 1 2 AOI21D0BWP7T $T=182960 200320 0 180 $X=179870 $Y=196110
X884 857 858 860 271 1 2 AOI21D0BWP7T $T=225520 168960 0 0 $X=225230 $Y=168725
X885 865 864 274 863 1 2 AOI21D0BWP7T $T=231680 184640 1 180 $X=228590 $Y=184405
X886 278 275 276 862 1 2 AOI21D0BWP7T $T=232800 200320 0 180 $X=229710 $Y=196110
X887 866 869 284 872 1 2 AOI21D0BWP7T $T=234480 192480 0 0 $X=234190 $Y=192245
X888 875 888 316 325 1 2 AOI21D0BWP7T $T=280400 184640 0 0 $X=280110 $Y=184405
X889 780 83 95 39 2 1 41 NR4D1BWP7T $T=85520 176800 1 180 $X=79630 $Y=176565
X890 790 125 16 792 2 1 19 NR4D1BWP7T $T=100080 192480 1 0 $X=99790 $Y=188270
X891 72 113 127 784 2 1 143 NR4D1BWP7T $T=105120 184640 0 0 $X=104830 $Y=184405
X892 144 83 142 794 2 1 118 NR4D1BWP7T $T=107920 176800 1 0 $X=107630 $Y=172590
X893 153 143 766 777 2 1 798 NR4D1BWP7T $T=121920 192480 1 0 $X=121630 $Y=188270
X894 804 122 82 177 2 1 799 NR4D1BWP7T $T=135360 184640 1 0 $X=135070 $Y=180430
X895 65 49 61 2 1 769 AN3D1BWP7T $T=59200 192480 1 180 $X=55550 $Y=192245
X896 762 767 68 2 1 71 AN3D1BWP7T $T=58080 192480 1 0 $X=57790 $Y=188270
X897 760 82 36 83 2 1 87 OR4D1BWP7T $T=67600 200320 1 0 $X=67310 $Y=196110
X898 69 88 83 94 2 1 782 OR4D1BWP7T $T=79920 200320 1 0 $X=79630 $Y=196110
X899 3 2 14 17 23 1 AOI21D2BWP7T $T=21120 176800 1 0 $X=20830 $Y=172590
X900 766 2 35 34 4 1 AOI21D2BWP7T $T=42960 184640 0 180 $X=37630 $Y=180430
X901 768 2 800 174 54 1 AOI21D2BWP7T $T=134240 176800 1 0 $X=133950 $Y=172590
X902 4 1 7 9 2 ND2D1BWP7T $T=21680 184640 1 0 $X=21390 $Y=180430
X903 5 1 11 15 2 ND2D1BWP7T $T=22240 192480 0 0 $X=21950 $Y=192245
X904 758 1 26 15 2 ND2D1BWP7T $T=29520 168960 1 180 $X=26990 $Y=168725
X905 24 1 21 23 2 ND2D1BWP7T $T=30080 184640 0 180 $X=27550 $Y=180430
X906 24 1 18 28 2 ND2D1BWP7T $T=27840 184640 0 0 $X=27550 $Y=184405
X907 23 1 761 31 2 ND2D1BWP7T $T=28960 176800 1 0 $X=28670 $Y=172590
X908 4 1 30 17 2 ND2D1BWP7T $T=28960 176800 0 0 $X=28670 $Y=176565
X909 38 1 764 17 2 ND2D1BWP7T $T=41840 176800 1 180 $X=39310 $Y=176565
X910 4 1 37 31 2 ND2D1BWP7T $T=40160 176800 1 0 $X=39870 $Y=172590
X911 767 1 39 7 2 ND2D1BWP7T $T=43520 184640 1 180 $X=40990 $Y=184405
X912 764 1 41 37 2 ND2D1BWP7T $T=42400 176800 1 0 $X=42110 $Y=172590
X913 4 1 44 5 2 ND2D1BWP7T $T=42960 192480 0 0 $X=42670 $Y=192245
X914 4 1 43 46 2 ND2D1BWP7T $T=43520 184640 0 0 $X=43230 $Y=184405
X915 764 1 53 43 2 ND2D1BWP7T $T=46320 200320 1 0 $X=46030 $Y=196110
X916 4 1 49 758 2 ND2D1BWP7T $T=46880 168960 0 0 $X=46590 $Y=168725
X917 34 1 50 52 2 ND2D1BWP7T $T=46880 184640 1 0 $X=46590 $Y=180430
X918 24 1 56 52 2 ND2D1BWP7T $T=49680 184640 1 0 $X=49390 $Y=180430
X919 52 1 63 46 2 ND2D1BWP7T $T=53040 184640 1 0 $X=52750 $Y=180430
X920 28 1 767 31 2 ND2D1BWP7T $T=56960 176800 0 180 $X=54430 $Y=172590
X921 38 1 64 46 2 ND2D1BWP7T $T=55840 176800 0 0 $X=55550 $Y=176565
X922 758 1 67 23 2 ND2D1BWP7T $T=57520 176800 1 0 $X=57230 $Y=172590
X923 29 1 66 761 2 ND2D1BWP7T $T=57520 184640 1 0 $X=57230 $Y=180430
X924 28 1 65 46 2 ND2D1BWP7T $T=60320 168960 1 180 $X=57790 $Y=168725
X925 34 1 75 23 2 ND2D1BWP7T $T=58640 176800 0 0 $X=58350 $Y=176565
X926 54 1 29 77 2 ND2D1BWP7T $T=61440 184640 1 0 $X=61150 $Y=180430
X927 758 1 68 28 2 ND2D1BWP7T $T=63120 176800 1 0 $X=62830 $Y=172590
X928 24 1 776 15 2 ND2D1BWP7T $T=68160 176800 1 0 $X=67870 $Y=172590
X929 54 1 81 46 2 ND2D1BWP7T $T=70400 184640 0 180 $X=67870 $Y=180430
X930 54 1 12 758 2 ND2D1BWP7T $T=69280 176800 0 0 $X=68990 $Y=176565
X931 31 1 85 15 2 ND2D1BWP7T $T=72640 168960 1 180 $X=70110 $Y=168725
X932 34 1 773 15 2 ND2D1BWP7T $T=73200 176800 0 180 $X=70670 $Y=172590
X933 54 1 778 31 2 ND2D1BWP7T $T=82720 176800 1 0 $X=82430 $Y=172590
X934 758 1 101 38 2 ND2D1BWP7T $T=86080 176800 0 0 $X=85790 $Y=176565
X935 778 1 784 65 2 ND2D1BWP7T $T=92240 184640 0 0 $X=91950 $Y=184405
X936 54 1 102 24 2 ND2D1BWP7T $T=98960 176800 0 180 $X=96430 $Y=172590
X937 758 1 788 132 2 ND2D1BWP7T $T=102880 176800 0 0 $X=102590 $Y=176565
X938 24 1 84 132 2 ND2D1BWP7T $T=107360 176800 1 180 $X=104830 $Y=176565
X939 788 1 133 134 2 ND2D1BWP7T $T=105120 200320 1 0 $X=104830 $Y=196110
X940 132 1 58 31 2 ND2D1BWP7T $T=106240 168960 0 0 $X=105950 $Y=168725
X941 137 1 774 141 2 ND2D1BWP7T $T=108480 168960 0 0 $X=108190 $Y=168725
X942 58 1 798 796 2 ND2D1BWP7T $T=122480 176800 0 0 $X=122190 $Y=176565
X943 217 1 222 194 2 ND2D1BWP7T $T=169520 176800 1 0 $X=169230 $Y=172590
X944 227 1 223 205 2 ND2D1BWP7T $T=174000 168960 0 0 $X=173710 $Y=168725
X945 205 1 824 806 2 ND2D1BWP7T $T=177360 176800 0 0 $X=177070 $Y=176565
X946 200 1 825 221 2 ND2D1BWP7T $T=179600 192480 0 0 $X=179310 $Y=192245
X947 206 1 834 221 2 ND2D1BWP7T $T=191360 192480 0 180 $X=188830 $Y=188270
X948 250 1 843 806 2 ND2D1BWP7T $T=199200 184640 1 180 $X=196670 $Y=184405
X949 187 1 251 831 2 ND2D1BWP7T $T=208160 192480 0 180 $X=205630 $Y=188270
X950 831 1 845 194 2 ND2D1BWP7T $T=208720 184640 1 0 $X=208430 $Y=180430
X951 846 1 262 263 2 ND2D1BWP7T $T=215440 184640 1 0 $X=215150 $Y=180430
X952 102 1 58 145 2 794 149 OAI211D1BWP7T $T=110720 168960 0 0 $X=110430 $Y=168725
X953 79 1 91 129 2 799 109 OAI211D1BWP7T $T=123600 176800 1 0 $X=123310 $Y=172590
X954 813 1 809 201 2 203 187 OAI211D1BWP7T $T=156640 200320 0 180 $X=152990 $Y=196110
X955 826 1 828 205 2 242 219 OAI211D1BWP7T $T=185760 192480 0 0 $X=185470 $Y=192245
X956 843 1 834 235 2 840 207 OAI211D1BWP7T $T=196960 184640 1 180 $X=193310 $Y=184405
X957 845 1 812 178 2 846 258 OAI211D1BWP7T $T=208720 184640 0 0 $X=208430 $Y=184405
X958 845 1 812 178 2 851 258 OAI211D1BWP7T $T=217680 192480 1 0 $X=217390 $Y=188270
X959 845 1 812 178 2 267 258 OAI211D1BWP7T $T=218800 184640 0 0 $X=218510 $Y=184405
X960 262 1 853 855 2 854 268 OAI211D1BWP7T $T=221600 192480 1 0 $X=221310 $Y=188270
X961 868 1 867 861 2 273 265 OAI211D1BWP7T $T=233360 176800 0 180 $X=229710 $Y=172590
X962 873 1 285 283 2 282 265 OAI211D1BWP7T $T=237840 184640 0 180 $X=234190 $Y=180430
X963 21 1 18 7 13 10 2 ND4D1BWP7T $T=26720 184640 1 180 $X=22510 $Y=184405
X964 30 1 29 27 757 760 2 ND4D1BWP7T $T=31200 192480 1 180 $X=26990 $Y=192245
X965 49 1 37 47 761 768 2 ND4D1BWP7T $T=51360 176800 0 180 $X=47150 $Y=172590
X966 75 1 773 761 43 771 2 ND4D1BWP7T $T=68720 184640 1 180 $X=64510 $Y=184405
X967 774 1 776 84 86 777 2 ND4D1BWP7T $T=69280 192480 1 0 $X=68990 $Y=188270
X968 68 1 102 64 773 103 2 ND4D1BWP7T $T=89440 176800 0 180 $X=85230 $Y=172590
X969 42 113 167 793 172 1 2 OAI31D1BWP7T $T=132000 200320 1 0 $X=131710 $Y=196110
X970 214 227 821 235 818 1 2 OAI31D1BWP7T $T=181840 176800 0 180 $X=177630 $Y=172590
X971 788 1 85 78 2 117 ND3D0BWP7T $T=98960 200320 0 180 $X=95870 $Y=196110
X972 187 1 180 216 2 827 ND3D0BWP7T $T=188560 192480 0 180 $X=185470 $Y=188270
X973 8 1 2 115 766 786 83 NR4D0BWP7T $T=93920 192480 1 0 $X=93630 $Y=188270
X974 766 1 2 775 122 165 42 NR4D0BWP7T $T=127520 192480 0 0 $X=127230 $Y=192245
X975 839 1 2 832 814 835 231 NR4D0BWP7T $T=191920 184640 0 180 $X=188270 $Y=180430
X976 840 1 2 829 220 844 249 NR4D0BWP7T $T=194160 176800 0 0 $X=193870 $Y=176565
X977 113 124 2 128 1 NR2D2BWP7T $T=99520 200320 1 0 $X=99230 $Y=196110
X978 229 223 2 807 1 NR2D2BWP7T $T=176800 176800 1 180 $X=172590 $Y=176565
X979 223 186 2 231 1 NR2D2BWP7T $T=178480 168960 0 0 $X=178190 $Y=168725
X980 197 180 2 239 1 NR2D2BWP7T $T=181840 192480 0 0 $X=181550 $Y=192245
X981 136 40 84 131 2 1 791 AN4D1BWP7T $T=107360 192480 1 180 $X=103150 $Y=192245
X982 234 222 824 827 2 1 237 AN4D1BWP7T $T=178480 184640 1 0 $X=178190 $Y=180430
X983 187 217 224 180 817 2 1 AOI31D1BWP7T $T=173440 192480 1 180 $X=169230 $Y=192245
X984 68 1 21 761 67 770 2 ND4D0BWP7T $T=62560 184640 1 180 $X=58910 $Y=184405
X985 774 1 12 56 73 765 2 ND4D0BWP7T $T=64800 192480 0 180 $X=61150 $Y=188270
X986 93 1 92 778 86 779 2 ND4D0BWP7T $T=83280 192480 0 180 $X=79630 $Y=188270
X987 84 1 50 105 107 783 2 ND4D0BWP7T $T=86080 192480 0 0 $X=85790 $Y=192245
X988 93 1 108 781 27 112 2 ND4D0BWP7T $T=90000 192480 1 0 $X=89710 $Y=188270
X989 105 1 786 787 148 797 2 ND4D0BWP7T $T=110720 192480 1 0 $X=110430 $Y=188270
X990 791 1 795 130 139 151 2 ND4D0BWP7T $T=111840 200320 1 0 $X=111550 $Y=196110
X991 136 1 71 800 155 158 2 ND4D0BWP7T $T=123600 200320 1 0 $X=123310 $Y=196110
X992 102 1 767 128 800 164 2 ND4D0BWP7T $T=128640 184640 0 0 $X=128350 $Y=184405
X993 804 1 130 128 168 169 2 ND4D0BWP7T $T=134800 192480 1 180 $X=131150 $Y=192245
X994 827 1 841 837 836 245 2 ND4D0BWP7T $T=195840 192480 1 180 $X=192190 $Y=192245
X995 178 194 828 2 1 240 OA21D0BWP7T $T=190240 200320 0 180 $X=186590 $Y=196110
X996 763 1 36 765 32 2 NR3D1BWP7T $T=42400 200320 0 180 $X=37630 $Y=196110
X997 195 1 180 189 191 2 NR3D1BWP7T $T=154400 192480 0 180 $X=149630 $Y=188270
X998 74 1 72 70 69 44 2 IND4D0BWP7T $T=63120 200320 0 180 $X=58910 $Y=196110
X999 143 1 89 139 793 126 2 IND4D0BWP7T $T=111280 200320 0 180 $X=107070 $Y=196110
X1000 98 1 96 780 90 63 2 IND4D1BWP7T $T=86640 184640 0 180 $X=81870 $Y=180430
X1001 785 1 781 76 111 778 2 IND4D1BWP7T $T=96720 176800 0 180 $X=91950 $Y=172590
X1002 798 1 168 73 805 790 2 IND4D1BWP7T $T=130880 192480 1 0 $X=130590 $Y=188270
X1003 62 2 20 8 759 1 40 NR4D3BWP7T $T=55280 192480 0 180 $X=39310 $Y=188270
X1004 773 766 1 100 781 2 INR3D1BWP7T $T=84960 184640 0 0 $X=84670 $Y=184405
X1005 171 2 113 1 145 NR2XD1BWP7T $T=136480 176800 1 180 $X=132270 $Y=176565
X1006 178 2 246 1 192 NR2XD1BWP7T $T=198080 168960 1 180 $X=193870 $Y=168725
X1007 42 1 45 37 2 IND2D1BWP7T $T=43520 176800 0 0 $X=43230 $Y=176565
X1008 88 1 82 762 2 IND2D1BWP7T $T=73200 184640 0 180 $X=70110 $Y=180430
X1009 24 15 19 6 8 1 2 AO211D2BWP7T $T=27280 192480 0 180 $X=21950 $Y=188270
X1010 79 1 91 129 2 109 789 OAI211D0BWP7T $T=106240 168960 1 180 $X=102590 $Y=168725
X1011 79 1 91 129 2 109 803 OAI211D0BWP7T $T=127520 176800 1 0 $X=127230 $Y=172590
X1012 206 1 205 187 2 214 836 OAI211D0BWP7T $T=189120 192480 0 0 $X=188830 $Y=192245
X1013 843 1 842 235 2 214 248 OAI211D0BWP7T $T=199200 192480 1 180 $X=195550 $Y=192245
X1014 251 1 252 182 2 201 255 OAI211D0BWP7T $T=205920 200320 1 0 $X=205630 $Y=196110
X1015 824 1 826 229 232 234 2 OAI211D2BWP7T $T=182400 192480 0 180 $X=175950 $Y=188270
X1016 845 1 812 258 850 178 2 OAI211D2BWP7T $T=212080 184640 0 0 $X=211790 $Y=184405
X1017 195 193 817 814 1 2 208 AO211D0BWP7T $T=168400 192480 0 180 $X=164190 $Y=188270
X1018 200 202 807 815 1 2 225 AO211D0BWP7T $T=168400 192480 1 0 $X=168110 $Y=188270
X1019 254 2 831 259 194 189 1 AOI211D2BWP7T $T=207040 168960 0 0 $X=206750 $Y=168725
X1020 166 2 766 170 1 NR2D3BWP7T $T=130320 168960 0 0 $X=130030 $Y=168725
X1021 190 2 196 197 1 NR2D3BWP7T $T=148240 200320 1 0 $X=147950 $Y=196110
X1022 206 2 193 180 1 NR2D3BWP7T $T=168960 192480 1 180 $X=163630 $Y=192245
X1023 219 2 220 187 1 NR2D3BWP7T $T=169520 184640 0 0 $X=169230 $Y=184405
X1024 209 2 226 228 1 NR2D3BWP7T $T=179040 200320 0 180 $X=173710 $Y=196110
X1025 28 79 9 1 2 ND2D2BWP7T $T=64240 168960 0 0 $X=63950 $Y=168725
X1026 157 170 174 1 2 ND2D2BWP7T $T=141520 168960 1 180 $X=137310 $Y=168725
X1027 180 178 806 1 2 ND2D2BWP7T $T=144320 184640 1 180 $X=140110 $Y=184405
X1028 186 189 184 1 2 ND2D2BWP7T $T=146000 168960 0 0 $X=145710 $Y=168725
X1029 200 207 206 1 2 ND2D2BWP7T $T=167840 184640 1 180 $X=163630 $Y=184405
X1030 209 211 214 1 2 ND2D2BWP7T $T=167280 184640 1 0 $X=166990 $Y=180430
X1031 217 219 200 1 2 ND2D2BWP7T $T=171200 184640 1 0 $X=170910 $Y=180430
X1032 337 2 351 319 338 1 893 346 AOI221D1BWP7T $T=307280 168960 1 180 $X=301950 $Y=168725
X1033 333 2 419 413 412 1 425 427 AOI221D1BWP7T $T=375040 168960 0 0 $X=374750 $Y=168725
X1034 333 2 911 416 423 1 910 909 AOI221D1BWP7T $T=381200 176800 1 180 $X=375870 $Y=176565
X1035 333 2 442 452 451 1 446 914 AOI221D1BWP7T $T=396880 184640 0 0 $X=396590 $Y=184405
X1036 16 1 2 775 106 104 NR3D0BWP7T $T=86080 200320 1 0 $X=85790 $Y=196110
X1037 62 1 2 118 100 787 NR3D0BWP7T $T=95600 184640 0 0 $X=95310 $Y=184405
X1038 150 1 2 114 122 795 NR3D0BWP7T $T=115200 192480 1 180 $X=112110 $Y=192245
X1039 17 23 1 25 757 2 AOI21D1BWP7T $T=25040 176800 0 0 $X=24750 $Y=176565
X1040 216 217 1 180 830 2 AOI21D1BWP7T $T=185200 176800 0 0 $X=184910 $Y=176565
X1041 240 843 251 825 260 1 2 ND4D2BWP7T $T=209840 200320 1 0 $X=209550 $Y=196110
X1042 27 1 792 33 156 157 2 OAI31D2BWP7T $T=128640 184640 1 180 $X=121630 $Y=184405
X1043 764 1 55 769 2 60 ND3D1BWP7T $T=49680 192480 0 0 $X=49390 $Y=192245
X1044 772 1 97 781 2 99 ND3D1BWP7T $T=83280 192480 1 0 $X=82990 $Y=188270
X1045 121 2 147 146 1 796 24 AOI211D1BWP7T $T=114640 184640 0 180 $X=110990 $Y=180430
X1046 802 2 60 175 1 176 801 AOI211D1BWP7T $T=135360 192480 1 0 $X=135070 $Y=188270
X1047 215 2 819 182 1 818 200 AOI211D1BWP7T $T=167840 168960 0 0 $X=167550 $Y=168725
X1048 869 2 864 865 1 853 277 AOI211D1BWP7T $T=235600 192480 0 180 $X=231950 $Y=188270
X1049 287 2 870 281 1 867 279 AOI211D1BWP7T $T=237280 168960 1 180 $X=233630 $Y=168725
X1050 67 2 78 25 1 INR2D1BWP7T $T=64240 192480 0 0 $X=63950 $Y=192245
X1051 186 239 806 241 243 1 2 244 AO221D0BWP7T $T=185200 168960 0 0 $X=184910 $Y=168725
X1052 295 296 300 878 2 1 297 DFCND1BWP7T $T=250720 192480 1 0 $X=250430 $Y=188270
X1053 45 1 2 66 77 772 80 AOI211XD0BWP7T $T=63680 176800 0 0 $X=63390 $Y=176565
X1054 121 1 2 784 5 110 38 AOI211XD0BWP7T $T=97280 184640 0 180 $X=93630 $Y=180430
X1055 771 1 2 121 150 154 156 AOI211XD0BWP7T $T=121920 184640 1 0 $X=121630 $Y=180430
X1056 181 1 2 807 182 809 806 AOI211XD0BWP7T $T=142640 192480 1 0 $X=142350 $Y=188270
X1057 821 1 2 231 205 820 209 AOI211XD0BWP7T $T=177920 176800 0 180 $X=174270 $Y=172590
X1058 443 912 393 444 441 1 2 DFCND2BWP7T $T=404160 176800 1 180 $X=389310 $Y=176565
X1059 443 457 393 448 445 1 2 DFCND2BWP7T $T=405840 192480 0 180 $X=390990 $Y=188270
X1060 85 1 98 33 109 2 OAI21D2BWP7T $T=87760 168960 0 0 $X=87470 $Y=168725
X1061 767 1 121 160 159 2 OAI21D2BWP7T $T=130320 184640 0 180 $X=124990 $Y=180430
X1062 371 1 366 367 898 2 OAI21D2BWP7T $T=319600 192480 0 180 $X=314270 $Y=188270
X1063 902 1 386 367 901 2 OAI21D2BWP7T $T=342560 184640 1 180 $X=337230 $Y=184405
X1064 915 1 460 367 465 2 OAI21D2BWP7T $T=408640 192480 1 180 $X=403310 $Y=192245
X1065 464 276 1 461 456 2 IOA21D1BWP7T $T=405840 168960 1 180 $X=402190 $Y=168725
X1066 201 192 1 211 2 815 195 OAI22D1BWP7T $T=163920 200320 1 0 $X=163630 $Y=196110
X1067 226 205 1 222 2 829 180 OAI22D1BWP7T $T=181280 176800 0 0 $X=180990 $Y=176565
X1068 806 234 1 197 2 832 217 OAI22D1BWP7T $T=188560 184640 0 180 $X=184350 $Y=180430
X1069 247 178 1 201 2 839 187 OAI22D1BWP7T $T=196960 192480 0 180 $X=192750 $Y=188270
X1070 852 265 1 271 2 862 859 OAI22D1BWP7T $T=226640 184640 1 0 $X=226350 $Y=180430
X1071 889 265 1 325 2 880 887 OAI22D1BWP7T $T=282080 168960 1 180 $X=277870 $Y=168725
X1072 322 332 320 891 337 1 2 341 AO221D1BWP7T $T=291600 192480 0 0 $X=291310 $Y=192245
X1073 331 856 334 894 333 1 2 350 AO221D1BWP7T $T=300560 176800 1 0 $X=300270 $Y=172590
X1074 361 364 365 897 333 1 2 370 AO221D1BWP7T $T=312320 200320 1 0 $X=312030 $Y=196110
X1075 368 860 896 899 337 1 2 378 AO221D1BWP7T $T=316800 176800 1 0 $X=316510 $Y=172590
X1076 387 389 388 391 333 1 2 392 AO221D1BWP7T $T=337520 192480 0 0 $X=337230 $Y=192245
X1077 421 424 422 426 428 1 2 430 AO221D1BWP7T $T=375600 192480 0 0 $X=375310 $Y=192245
X1078 496 501 917 921 333 1 2 505 AO221D1BWP7T $T=438320 200320 1 0 $X=438030 $Y=196110
X1079 509 486 923 924 333 1 2 513 AO221D1BWP7T $T=445600 192480 1 0 $X=445310 $Y=188270
X1080 515 516 517 925 428 1 2 526 AO221D1BWP7T $T=459040 200320 1 0 $X=458750 $Y=196110
X1081 295 303 300 294 2 1 292 DFCND0BWP7T $T=262480 184640 0 180 $X=249310 $Y=180430
X1082 295 305 300 291 2 1 874 DFCND0BWP7T $T=264160 192480 1 180 $X=250990 $Y=192245
X1083 295 883 300 879 2 1 877 DFCND0BWP7T $T=272560 176800 1 180 $X=259390 $Y=176565
X1084 295 881 300 313 2 1 885 DFCND0BWP7T $T=264160 184640 0 0 $X=263870 $Y=184405
X1085 400 905 393 402 2 1 394 DFCND0BWP7T $T=364400 176800 0 180 $X=351230 $Y=172590
X1086 443 447 393 913 2 1 458 DFCND0BWP7T $T=390720 200320 1 0 $X=390430 $Y=196110
X1087 886 315 182 314 308 313 2 882 1 OA222D0BWP7T $T=275360 192480 1 180 $X=268910 $Y=192245
X1088 321 315 182 318 309 310 2 884 1 OA222D0BWP7T $T=277600 176800 0 180 $X=271150 $Y=172590
X1089 770 2 39 1 51 5 54 AOI211XD1BWP7T $T=54720 184640 1 180 $X=47710 $Y=184405
X1090 188 2 807 1 198 194 189 AOI211XD1BWP7T $T=146560 184640 1 0 $X=146270 $Y=180430
X1091 880 2 870 1 307 279 298 AOI211XD1BWP7T $T=259680 176800 1 0 $X=259390 $Y=172590
X1092 315 317 1 301 311 308 291 2 304 OAI222D2BWP7T $T=274800 200320 0 180 $X=264430 $Y=196110
X1093 315 319 1 182 312 309 878 2 306 OAI222D2BWP7T $T=276480 168960 1 180 $X=266110 $Y=168725
X1094 180 204 206 1 2 ND2D1P5BWP7T $T=163920 168960 0 0 $X=163630 $Y=168725
X1095 99 2 122 801 1 173 157 AOI211XD2BWP7T $T=134800 192480 0 0 $X=134510 $Y=192245
X1096 810 2 811 193 1 812 202 AOI211XD2BWP7T $T=144320 184640 0 0 $X=144030 $Y=184405
X1097 1 2 ICV_23 $T=119120 192480 0 0 $X=118830 $Y=192245
X1098 1 2 ICV_23 $T=195280 200320 1 0 $X=194990 $Y=196110
X1099 1 2 ICV_23 $T=203120 176800 0 0 $X=202830 $Y=176565
X1100 1 2 ICV_23 $T=245120 168960 0 0 $X=244830 $Y=168725
X1101 1 2 ICV_23 $T=245120 200320 1 0 $X=244830 $Y=196110
X1102 1 2 ICV_23 $T=277600 176800 1 0 $X=277310 $Y=172590
X1103 1 2 ICV_23 $T=293840 176800 1 0 $X=293550 $Y=172590
X1104 1 2 ICV_23 $T=293840 176800 0 0 $X=293550 $Y=176565
X1105 1 2 ICV_23 $T=296640 184640 0 0 $X=296350 $Y=184405
X1106 1 2 ICV_23 $T=296640 192480 1 0 $X=296350 $Y=188270
X1107 1 2 ICV_23 $T=329120 184640 0 0 $X=328830 $Y=184405
X1108 1 2 ICV_23 $T=329120 192480 0 0 $X=328830 $Y=192245
X1109 1 2 ICV_23 $T=342560 184640 0 0 $X=342270 $Y=184405
X1110 1 2 ICV_23 $T=353760 184640 0 0 $X=353470 $Y=184405
X1111 1 2 ICV_23 $T=362160 192480 1 0 $X=361870 $Y=188270
X1112 1 2 ICV_23 $T=371120 192480 1 0 $X=370830 $Y=188270
X1113 1 2 ICV_23 $T=388480 168960 0 0 $X=388190 $Y=168725
X1114 1 2 ICV_23 $T=404160 176800 0 0 $X=403870 $Y=176565
X1115 1 2 ICV_23 $T=413120 168960 0 0 $X=412830 $Y=168725
X1116 1 2 ICV_23 $T=413120 176800 0 0 $X=412830 $Y=176565
X1117 1 2 ICV_23 $T=413120 184640 1 0 $X=412830 $Y=180430
X1118 1 2 ICV_23 $T=413120 200320 1 0 $X=412830 $Y=196110
X1119 1 2 ICV_23 $T=426560 200320 1 0 $X=426270 $Y=196110
X1120 1 2 ICV_23 $T=427680 176800 0 0 $X=427390 $Y=176565
X1121 1 2 ICV_23 $T=429920 168960 0 0 $X=429630 $Y=168725
X1122 1 2 ICV_23 $T=442800 192480 0 0 $X=442510 $Y=192245
X1123 1 2 ICV_23 $T=446160 168960 0 0 $X=445870 $Y=168725
X1124 1 2 ICV_23 $T=446160 200320 1 0 $X=445870 $Y=196110
X1125 1 2 ICV_23 $T=447280 176800 1 0 $X=446990 $Y=172590
X1126 403 1 263 404 2 CKND2D2BWP7T $T=354880 184640 0 180 $X=350670 $Y=180430
X1127 328 329 886 890 333 336 1 2 AO221D2BWP7T $T=289920 184640 0 0 $X=289630 $Y=184405
X1128 339 274 335 895 333 355 1 2 AO221D2BWP7T $T=303360 184640 0 0 $X=303070 $Y=184405
X1129 479 503 922 508 333 512 1 2 AO221D2BWP7T $T=440560 176800 1 0 $X=440270 $Y=172590
X1130 192 1 184 185 187 178 2 OAI22D2BWP7T $T=152720 176800 0 180 $X=145710 $Y=172590
X1131 381 367 1 2 CKND8BWP7T $T=347600 168960 1 180 $X=340590 $Y=168725
X1132 333 2 499 1 507 NR2XD3BWP7T $T=446160 168960 1 180 $X=437470 $Y=168725
X1133 428 2 520 1 523 NR2D5BWP7T $T=470800 168960 1 180 $X=462110 $Y=168725
X1134 428 2 519 1 524 NR2D5BWP7T $T=470800 176800 0 180 $X=462110 $Y=172590
X1135 428 2 521 1 525 NR2D5BWP7T $T=470800 192480 0 180 $X=462110 $Y=188270
X1136 428 522 514 1 2 INR2XD4BWP7T $T=470800 176800 1 180 $X=457630 $Y=176565
X1137 197 1 256 2 849 OR2D1BWP7T $T=218240 184640 1 0 $X=217950 $Y=180430
X1138 317 1 333 2 340 OR2D1BWP7T $T=294400 184640 1 0 $X=294110 $Y=180430
.ENDS
***************************************
.SUBCKT ICV_31 1 2
** N=2 EP=2 IP=4 FDC=2
X1 2 1 DCAPBWP7T $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ND2D3BWP7T A2 VSS ZN A1 VDD
** N=6 EP=5 IP=0 FDC=12
M0 6 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=620 $Y=345 $D=0
M1 VSS A2 6 VSS N L=1.8e-07 W=1e-06 $X=1340 $Y=345 $D=0
M2 6 A2 VSS VSS N L=1.8e-07 W=1e-06 $X=2060 $Y=345 $D=0
M3 ZN A1 6 VSS N L=1.8e-07 W=1e-06 $X=2780 $Y=345 $D=0
M4 6 A1 ZN VSS N L=1.8e-07 W=1e-06 $X=3500 $Y=345 $D=0
M5 ZN A1 6 VSS N L=1.8e-07 W=1e-06 $X=4220 $Y=345 $D=0
M6 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=620 $Y=2205 $D=16
M7 VDD A2 ZN VDD P L=1.8e-07 W=1.37e-06 $X=1340 $Y=2205 $D=16
M8 ZN A2 VDD VDD P L=1.8e-07 W=1.37e-06 $X=2060 $Y=2205 $D=16
M9 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=2780 $Y=2205 $D=16
M10 ZN A1 VDD VDD P L=1.8e-07 W=1.37e-06 $X=3500 $Y=2205 $D=16
M11 VDD A1 ZN VDD P L=1.8e-07 W=1.37e-06 $X=4220 $Y=2205 $D=16
.ENDS
***************************************
.SUBCKT ICV_32 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480
+ 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500
+ 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520
+ 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540
+ 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560
+ 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580
+ 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600
+ 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620
+ 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640
+ 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660
+ 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680
+ 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700
+ 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720
+ 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740
+ 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760
+ 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780
+ 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800
+ 801
** N=1410 EP=801 IP=6557 FDC=10406
M0 918 28 919 1 N L=1.8e-07 W=1e-06 $X=26995 $Y=128415 $D=0
M1 919 31 918 1 N L=1.8e-07 W=1e-06 $X=27715 $Y=128415 $D=0
M2 1 925 919 1 N L=1.8e-07 W=1e-06 $X=28435 $Y=128415 $D=0
M3 1391 35 1 1 N L=1.8e-07 W=1e-06 $X=29195 $Y=128415 $D=0
M4 925 23 1391 1 N L=1.8e-07 W=1e-06 $X=29755 $Y=128415 $D=0
M5 1010 185 1 1 N L=1.8e-07 W=1e-06 $X=86185 $Y=122265 $D=0
M6 1 980 1010 1 N L=1.8e-07 W=1e-06 $X=86905 $Y=122265 $D=0
M7 1010 999 1 1 N L=1.8e-07 W=1e-06 $X=87705 $Y=122265 $D=0
M8 1 181 1010 1 N L=1.8e-07 W=1e-06 $X=88425 $Y=122265 $D=0
M9 193 1010 1 1 N L=1.8e-07 W=1e-06 $X=91520 $Y=122265 $D=0
M10 1 1010 193 1 N L=1.8e-07 W=1e-06 $X=92240 $Y=122265 $D=0
M11 193 1010 1 1 N L=1.8e-07 W=1e-06 $X=92960 $Y=122265 $D=0
M12 1 1010 193 1 N L=1.8e-07 W=1e-06 $X=93680 $Y=122265 $D=0
M13 417 359 1157 1 N L=1.8e-07 W=1e-06 $X=187575 $Y=144095 $D=0
M14 1157 359 417 1 N L=1.8e-07 W=1e-06 $X=188295 $Y=144095 $D=0
M15 417 359 1157 1 N L=1.8e-07 W=1e-06 $X=189015 $Y=144095 $D=0
M16 1157 359 417 1 N L=1.8e-07 W=1e-06 $X=189735 $Y=144095 $D=0
M17 417 359 1157 1 N L=1.8e-07 W=1e-06 $X=190455 $Y=144095 $D=0
M18 1157 359 417 1 N L=1.8e-07 W=1e-06 $X=191175 $Y=144095 $D=0
M19 417 359 1157 1 N L=1.8e-07 W=1e-06 $X=191895 $Y=144095 $D=0
M20 1157 359 417 1 N L=1.8e-07 W=1e-06 $X=192620 $Y=144095 $D=0
M21 1 388 1157 1 N L=1.8e-07 W=1e-06 $X=193340 $Y=144095 $D=0
M22 1157 388 1 1 N L=1.8e-07 W=1e-06 $X=194060 $Y=144095 $D=0
M23 1 388 1157 1 N L=1.8e-07 W=1e-06 $X=194780 $Y=144095 $D=0
M24 1157 388 1 1 N L=1.8e-07 W=1e-06 $X=195500 $Y=144095 $D=0
M25 1 388 1157 1 N L=1.8e-07 W=1e-06 $X=196220 $Y=144095 $D=0
M26 1157 388 1 1 N L=1.8e-07 W=1e-06 $X=196940 $Y=144095 $D=0
M27 1 388 1157 1 N L=1.8e-07 W=1e-06 $X=197660 $Y=144095 $D=0
M28 1157 388 1 1 N L=1.8e-07 W=1e-06 $X=198380 $Y=144095 $D=0
M29 1 355 1164 1 N L=1.8e-07 W=5e-07 $X=208220 $Y=122425 $D=0
M30 1392 388 1 1 N L=1.8e-07 W=5.7e-07 $X=208980 $Y=122695 $D=0
M31 1169 355 1392 1 N L=1.8e-07 W=5.7e-07 $X=209410 $Y=122695 $D=0
M32 1393 1164 1169 1 N L=1.8e-07 W=4.2e-07 $X=210170 $Y=122570 $D=0
M33 1 1180 1393 1 N L=1.8e-07 W=4.2e-07 $X=210600 $Y=122570 $D=0
M34 1 374 1166 1 N L=1.8e-07 W=5e-07 $X=211860 $Y=122900 $D=0
M35 1167 1166 1 1 N L=1.8e-07 W=5e-07 $X=212465 $Y=122900 $D=0
M36 1172 1166 1169 1 N L=1.8e-07 W=7.4e-07 $X=213885 $Y=122495 $D=0
M37 1394 1167 1172 1 N L=1.8e-07 W=4.2e-07 $X=214715 $Y=122815 $D=0
M38 1395 382 1394 1 N L=1.8e-07 W=4.2e-07 $X=215175 $Y=122815 $D=0
M39 1 1176 1395 1 N L=1.8e-07 W=4.2e-07 $X=215635 $Y=122815 $D=0
M40 1176 1172 1 1 N L=1.8e-07 W=5.4e-07 $X=216495 $Y=122695 $D=0
M41 1182 1167 1176 1 N L=1.8e-07 W=9.1e-07 $X=217370 $Y=122325 $D=0
M42 1180 1166 1182 1 N L=1.8e-07 W=4.2e-07 $X=218135 $Y=122815 $D=0
M43 1 1188 1180 1 N L=1.8e-07 W=4.2e-07 $X=219925 $Y=122775 $D=0
M44 1396 382 1 1 N L=1.8e-07 W=9.3e-07 $X=220570 $Y=122265 $D=0
M45 1188 1182 1396 1 N L=1.8e-07 W=1e-06 $X=221210 $Y=122265 $D=0
M46 1 1180 1186 1 N L=1.8e-07 W=9.4e-07 $X=222880 $Y=122325 $D=0
M47 1181 1188 1 1 N L=1.8e-07 W=1e-06 $X=223600 $Y=122265 $D=0
M48 1268 484 1 1 N L=1.8e-07 W=5.7e-07 $X=300730 $Y=152365 $D=0
M49 1 1266 1268 1 N L=1.8e-07 W=5.7e-07 $X=301450 $Y=152365 $D=0
M50 557 1268 1 1 N L=1.8e-07 W=1e-06 $X=302230 $Y=151935 $D=0
M51 1 1262 557 1 N L=1.8e-07 W=1e-06 $X=302950 $Y=151935 $D=0
M52 1369 503 1367 1 N L=1.8e-07 W=1e-06 $X=398060 $Y=137945 $D=0
M53 1367 692 1369 1 N L=1.8e-07 W=1e-06 $X=398780 $Y=137945 $D=0
M54 1367 1356 1371 1 N L=1.8e-07 W=1e-06 $X=400080 $Y=137945 $D=0
M55 1371 526 1367 1 N L=1.8e-07 W=1e-06 $X=400800 $Y=137945 $D=0
M56 1 640 1371 1 N L=1.8e-07 W=1e-06 $X=401520 $Y=137945 $D=0
M57 1371 698 1 1 N L=1.8e-07 W=1e-06 $X=402240 $Y=137945 $D=0
M58 1397 28 2 2 P L=1.8e-07 W=1.37e-06 $X=26875 $Y=126185 $D=16
M59 918 31 1397 2 P L=1.8e-07 W=1.37e-06 $X=27475 $Y=126185 $D=16
M60 2 925 918 2 P L=1.8e-07 W=1.37e-06 $X=28195 $Y=126185 $D=16
M61 925 35 2 2 P L=1.8e-07 W=1.37e-06 $X=29035 $Y=126185 $D=16
M62 2 23 925 2 P L=1.8e-07 W=1.37e-06 $X=29755 $Y=126185 $D=16
M63 1398 185 2 2 P L=1.8e-07 W=1.37e-06 $X=86245 $Y=124125 $D=16
M64 1399 980 1398 2 P L=1.8e-07 W=1.37e-06 $X=86845 $Y=124125 $D=16
M65 1400 999 1399 2 P L=1.8e-07 W=1.37e-06 $X=87445 $Y=124125 $D=16
M66 1010 181 1400 2 P L=1.8e-07 W=1.37e-06 $X=88045 $Y=124125 $D=16
M67 1401 181 1010 2 P L=1.8e-07 W=1.37e-06 $X=88845 $Y=124125 $D=16
M68 1402 999 1401 2 P L=1.8e-07 W=1.37e-06 $X=89470 $Y=124125 $D=16
M69 1403 980 1402 2 P L=1.8e-07 W=1.37e-06 $X=90095 $Y=124125 $D=16
M70 2 185 1403 2 P L=1.8e-07 W=1.37e-06 $X=90720 $Y=124125 $D=16
M71 193 1010 2 2 P L=1.8e-07 W=1.37e-06 $X=91520 $Y=124125 $D=16
M72 2 1010 193 2 P L=1.8e-07 W=1.37e-06 $X=92240 $Y=124125 $D=16
M73 193 1010 2 2 P L=1.8e-07 W=1.37e-06 $X=92960 $Y=124125 $D=16
M74 2 1010 193 2 P L=1.8e-07 W=1.37e-06 $X=93680 $Y=124125 $D=16
M75 417 359 2 2 P L=1.8e-07 W=1.37e-06 $X=187575 $Y=141865 $D=16
M76 2 359 417 2 P L=1.8e-07 W=1.37e-06 $X=188295 $Y=141865 $D=16
M77 417 359 2 2 P L=1.8e-07 W=1.37e-06 $X=189015 $Y=141865 $D=16
M78 2 359 417 2 P L=1.8e-07 W=1.37e-06 $X=189735 $Y=141865 $D=16
M79 417 359 2 2 P L=1.8e-07 W=1.37e-06 $X=190455 $Y=141865 $D=16
M80 2 359 417 2 P L=1.8e-07 W=1.37e-06 $X=191175 $Y=141865 $D=16
M81 417 359 2 2 P L=1.8e-07 W=1.37e-06 $X=191895 $Y=141865 $D=16
M82 2 359 417 2 P L=1.8e-07 W=1.37e-06 $X=192620 $Y=141865 $D=16
M83 417 388 2 2 P L=1.8e-07 W=1.37e-06 $X=193340 $Y=141865 $D=16
M84 2 388 417 2 P L=1.8e-07 W=1.37e-06 $X=194060 $Y=141865 $D=16
M85 417 388 2 2 P L=1.8e-07 W=1.37e-06 $X=194780 $Y=141865 $D=16
M86 2 388 417 2 P L=1.8e-07 W=1.37e-06 $X=195500 $Y=141865 $D=16
M87 417 388 2 2 P L=1.8e-07 W=1.37e-06 $X=196220 $Y=141865 $D=16
M88 2 388 417 2 P L=1.8e-07 W=1.37e-06 $X=196940 $Y=141865 $D=16
M89 417 388 2 2 P L=1.8e-07 W=1.37e-06 $X=197660 $Y=141865 $D=16
M90 2 388 417 2 P L=1.8e-07 W=1.37e-06 $X=198380 $Y=141865 $D=16
M91 2 355 1164 2 P L=1.8e-07 W=6.85e-07 $X=208220 $Y=124750 $D=16
M92 1404 388 2 2 P L=1.8e-07 W=7.5e-07 $X=208980 $Y=124315 $D=16
M93 1169 1164 1404 2 P L=1.8e-07 W=7.5e-07 $X=209410 $Y=124315 $D=16
M94 1405 355 1169 2 P L=1.8e-07 W=4.2e-07 $X=210130 $Y=124645 $D=16
M95 2 1180 1405 2 P L=1.8e-07 W=4.2e-07 $X=210560 $Y=124645 $D=16
M96 2 374 1166 2 P L=1.8e-07 W=6.85e-07 $X=211860 $Y=124265 $D=16
M97 1167 1166 2 2 P L=1.8e-07 W=6.85e-07 $X=212470 $Y=124265 $D=16
M98 1172 1167 1169 2 P L=1.8e-07 W=7.8e-07 $X=213890 $Y=124265 $D=16
M99 1170 1166 1172 2 P L=1.8e-07 W=4.2e-07 $X=214745 $Y=124265 $D=16
M100 2 382 1170 2 P L=1.8e-07 W=4.2e-07 $X=215465 $Y=124265 $D=16
M101 1170 1176 2 2 P L=1.8e-07 W=4.2e-07 $X=216065 $Y=124265 $D=16
M102 1176 1172 2 2 P L=1.8e-07 W=6.2e-07 $X=217335 $Y=124095 $D=16
M103 1182 1166 1176 2 P L=1.8e-07 W=6.2e-07 $X=218135 $Y=124095 $D=16
M104 1180 1167 1182 2 P L=1.8e-07 W=4.2e-07 $X=219050 $Y=124130 $D=16
M105 2 1188 1180 2 P L=1.8e-07 W=6.85e-07 $X=219925 $Y=124130 $D=16
M106 1188 382 2 2 P L=1.8e-07 W=4.2e-07 $X=220810 $Y=124740 $D=16
M107 2 1182 1188 2 P L=1.8e-07 W=1.03e-06 $X=221580 $Y=124130 $D=16
M108 2 1180 1186 2 P L=1.8e-07 W=1.37e-06 $X=222880 $Y=124125 $D=16
M109 1181 1188 2 2 P L=1.8e-07 W=1.37e-06 $X=223600 $Y=124125 $D=16
M110 1406 484 1268 2 P L=1.8e-07 W=8.1e-07 $X=300730 $Y=149705 $D=16
M111 2 1266 1406 2 P L=1.8e-07 W=8.1e-07 $X=301330 $Y=149705 $D=16
M112 1407 1268 2 2 P L=1.8e-07 W=1.37e-06 $X=302230 $Y=149705 $D=16
M113 557 1262 1407 2 P L=1.8e-07 W=1.37e-06 $X=302830 $Y=149705 $D=16
M114 1408 503 1369 2 P L=1.8e-07 W=1.295e-06 $X=398060 $Y=139880 $D=16
M115 2 692 1408 2 P L=1.8e-07 W=1.25e-06 $X=398780 $Y=139925 $D=16
M116 1409 1356 2 2 P L=1.8e-07 W=1.25e-06 $X=400080 $Y=139925 $D=16
M117 1369 526 1409 2 P L=1.8e-07 W=1.37e-06 $X=400800 $Y=139805 $D=16
M118 1410 640 1369 2 P L=1.8e-07 W=1.37e-06 $X=401600 $Y=139805 $D=16
M119 2 698 1410 2 P L=1.8e-07 W=1.37e-06 $X=402240 $Y=139805 $D=16
X189 1 798 ANTENNABWP7T $T=471920 168960 0 180 $X=470510 $Y=164750
X190 1 564 ANTENNABWP7T $T=473040 168960 0 180 $X=471630 $Y=164750
X191 1 551 ANTENNABWP7T $T=474160 168960 0 180 $X=472750 $Y=164750
X292 934 1 2 936 CKBD1BWP7T $T=41280 153280 0 0 $X=40990 $Y=153045
X293 955 1 2 978 CKBD1BWP7T $T=67040 137600 1 0 $X=66750 $Y=133390
X294 148 1 2 986 CKBD1BWP7T $T=69280 137600 1 0 $X=68990 $Y=133390
X295 186 1 2 1006 CKBD1BWP7T $T=92240 137600 0 180 $X=89710 $Y=133390
X296 1100 1 2 322 CKBD1BWP7T $T=144880 168960 1 0 $X=144590 $Y=164750
X297 1142 1 2 406 CKBD1BWP7T $T=189680 114080 1 180 $X=187150 $Y=113845
X298 1150 1 2 418 CKBD1BWP7T $T=194160 129760 0 180 $X=191630 $Y=125550
X299 1152 1 2 424 CKBD1BWP7T $T=196400 121920 0 180 $X=193870 $Y=117710
X300 447 1 2 448 CKBD1BWP7T $T=217680 121920 1 0 $X=217390 $Y=117710
X301 451 1 2 1183 CKBD1BWP7T $T=219920 129760 0 0 $X=219630 $Y=129525
X302 1174 1 2 454 CKBD1BWP7T $T=219920 161120 0 0 $X=219630 $Y=160885
X303 1204 1 2 500 CKBD1BWP7T $T=249040 114080 0 0 $X=248750 $Y=113845
X304 1211 1 2 509 CKBD1BWP7T $T=256320 145440 0 180 $X=253790 $Y=141230
X305 1239 1 2 452 CKBD1BWP7T $T=272560 145440 0 0 $X=272270 $Y=145205
X306 1240 1 2 510 CKBD1BWP7T $T=275360 106240 0 0 $X=275070 $Y=106005
X307 1275 1 2 573 CKBD1BWP7T $T=310640 106240 0 0 $X=310350 $Y=106005
X308 584 1 2 560 CKBD1BWP7T $T=319040 161120 0 180 $X=316510 $Y=156910
X309 591 1 2 1293 CKBD1BWP7T $T=331920 153280 0 0 $X=331630 $Y=153045
X310 616 1 2 600 CKBD1BWP7T $T=343680 161120 0 180 $X=341150 $Y=156910
X311 1144 1 2 1321 CKBD1BWP7T $T=357680 114080 0 180 $X=355150 $Y=109870
X312 1318 1 2 626 CKBD1BWP7T $T=358240 121920 0 180 $X=355710 $Y=117710
X313 638 1 2 634 CKBD1BWP7T $T=359920 168960 0 180 $X=357390 $Y=164750
X314 1354 1 2 684 CKBD1BWP7T $T=391840 145440 0 0 $X=391550 $Y=145205
X315 670 1 2 708 CKBD1BWP7T $T=418160 161120 0 180 $X=415630 $Y=156910
X316 739 1 2 738 CKBD1BWP7T $T=434960 129760 1 180 $X=432430 $Y=129525
X317 710 1 2 744 CKBD1BWP7T $T=437760 137600 0 180 $X=435230 $Y=133390
X318 15 1 2 31 INVD0BWP7T $T=25600 121920 0 0 $X=25310 $Y=121685
X319 3 1 2 931 INVD0BWP7T $T=37920 145440 0 0 $X=37630 $Y=145205
X320 49 1 2 928 INVD0BWP7T $T=43520 137600 1 180 $X=41550 $Y=137365
X321 44 1 2 933 INVD0BWP7T $T=45200 137600 1 180 $X=43230 $Y=137365
X322 59 1 2 73 INVD0BWP7T $T=46880 114080 0 0 $X=46590 $Y=113845
X323 944 1 2 963 INVD0BWP7T $T=57520 137600 1 0 $X=57230 $Y=133390
X324 107 1 2 962 INVD0BWP7T $T=59200 145440 0 180 $X=57230 $Y=141230
X325 957 1 2 121 INVD0BWP7T $T=60320 114080 1 0 $X=60030 $Y=109870
X326 153 1 2 985 INVD0BWP7T $T=71520 153280 0 0 $X=71230 $Y=153045
X327 159 1 2 992 INVD0BWP7T $T=81600 145440 1 180 $X=79630 $Y=145205
X328 966 1 2 154 INVD0BWP7T $T=86640 114080 1 180 $X=84670 $Y=113845
X329 1026 1 2 1029 INVD0BWP7T $T=103440 137600 1 0 $X=103150 $Y=133390
X330 202 1 2 225 INVD0BWP7T $T=104000 106240 0 0 $X=103710 $Y=106005
X331 1023 1 2 1030 INVD0BWP7T $T=107360 161120 1 0 $X=107070 $Y=156910
X332 254 1 2 1045 INVD0BWP7T $T=113520 145440 1 0 $X=113230 $Y=141230
X333 259 1 2 1049 INVD0BWP7T $T=121920 106240 0 0 $X=121630 $Y=106005
X334 1035 1 2 1048 INVD0BWP7T $T=121920 145440 1 0 $X=121630 $Y=141230
X335 143 1 2 270 INVD0BWP7T $T=123040 153280 1 0 $X=122750 $Y=149070
X336 1071 1 2 1070 INVD0BWP7T $T=133120 121920 0 180 $X=131150 $Y=117710
X337 296 1 2 1039 INVD0BWP7T $T=135920 114080 0 180 $X=133950 $Y=109870
X338 1031 1 2 1082 INVD0BWP7T $T=135360 137600 0 0 $X=135070 $Y=137365
X339 1075 1 2 1085 INVD0BWP7T $T=137040 137600 0 0 $X=136750 $Y=137365
X340 309 1 2 1081 INVD0BWP7T $T=143200 129760 0 180 $X=141230 $Y=125550
X341 338 1 2 318 INVD0BWP7T $T=153840 114080 1 0 $X=153550 $Y=109870
X342 1120 1 2 1114 INVD0BWP7T $T=156640 129760 1 180 $X=154670 $Y=129525
X343 1121 1 2 1120 INVD0BWP7T $T=157200 121920 0 180 $X=155230 $Y=117710
X344 316 1 2 1123 INVD0BWP7T $T=164480 121920 1 0 $X=164190 $Y=117710
X345 354 1 2 356 INVD0BWP7T $T=165040 168960 1 0 $X=164750 $Y=164750
X346 436 1 2 1162 INVD0BWP7T $T=209280 121920 0 180 $X=207310 $Y=117710
X347 453 1 2 449 INVD0BWP7T $T=221600 106240 1 180 $X=219630 $Y=106005
X348 1156 1 2 1185 INVD0BWP7T $T=221040 137600 0 0 $X=220750 $Y=137365
X349 457 1 2 1175 INVD0BWP7T $T=224400 106240 1 180 $X=222430 $Y=106005
X350 473 1 2 1194 INVD0BWP7T $T=233360 161120 0 0 $X=233070 $Y=160885
X351 1208 1 2 1205 INVD0BWP7T $T=254080 137600 1 180 $X=252110 $Y=137365
X352 1213 1 2 1215 INVD0BWP7T $T=255760 114080 0 0 $X=255470 $Y=113845
X353 1227 1 2 1210 INVD0BWP7T $T=264720 137600 0 180 $X=262750 $Y=133390
X354 1220 1 2 1223 INVD0BWP7T $T=263600 114080 0 0 $X=263310 $Y=113845
X355 1236 1 2 1231 INVD0BWP7T $T=273680 129760 0 180 $X=271710 $Y=125550
X356 1246 1 2 1249 INVD0BWP7T $T=281520 129760 1 0 $X=281230 $Y=125550
X357 1250 1 2 1255 INVD0BWP7T $T=289920 145440 1 0 $X=289630 $Y=141230
X358 1259 1 2 1256 INVD0BWP7T $T=294960 114080 0 180 $X=292990 $Y=109870
X359 549 1 2 550 INVD0BWP7T $T=297760 137600 1 0 $X=297470 $Y=133390
X360 553 1 2 556 INVD0BWP7T $T=303920 168960 0 180 $X=301950 $Y=164750
X361 558 1 2 1267 INVD0BWP7T $T=305040 114080 0 180 $X=303070 $Y=109870
X362 560 1 2 1270 INVD0BWP7T $T=308400 137600 1 180 $X=306430 $Y=137365
X363 551 1 2 1272 INVD0BWP7T $T=308960 161120 0 180 $X=306990 $Y=156910
X364 572 1 2 1278 INVD0BWP7T $T=323520 106240 1 180 $X=321550 $Y=106005
X365 596 1 2 599 INVD0BWP7T $T=331920 137600 1 0 $X=331630 $Y=133390
X366 600 1 2 1294 INVD0BWP7T $T=335280 114080 0 180 $X=333310 $Y=109870
X367 591 1 2 1297 INVD0BWP7T $T=335840 145440 0 0 $X=335550 $Y=145205
X368 1306 1 2 1298 INVD0BWP7T $T=339200 145440 1 180 $X=337230 $Y=145205
X369 1191 1 2 1295 INVD0BWP7T $T=340880 145440 0 180 $X=338910 $Y=141230
X370 530 1 2 1299 INVD0BWP7T $T=345360 137600 0 180 $X=343390 $Y=133390
X371 1310 1 2 1306 INVD0BWP7T $T=348160 153280 1 180 $X=346190 $Y=153045
X372 609 1 2 1301 INVD0BWP7T $T=350960 161120 1 180 $X=348990 $Y=160885
X373 1305 1 2 1319 INVD0BWP7T $T=352640 145440 1 0 $X=352350 $Y=141230
X374 1317 1 2 1334 INVD0BWP7T $T=364400 121920 0 0 $X=364110 $Y=121685
X375 1325 1 2 654 INVD0BWP7T $T=373920 161120 0 0 $X=373630 $Y=160885
X376 649 1 2 660 INVD0BWP7T $T=378960 168960 0 180 $X=376990 $Y=164750
X377 1341 1 2 1348 INVD0BWP7T $T=385120 129760 1 0 $X=384830 $Y=125550
X378 1359 1 2 1358 INVD0BWP7T $T=396880 137600 1 180 $X=394910 $Y=137365
X379 1363 1 2 691 INVD0BWP7T $T=399120 161120 1 180 $X=397150 $Y=160885
X380 702 1 2 1360 INVD0BWP7T $T=404720 106240 1 180 $X=402750 $Y=106005
X381 1369 1 2 1359 INVD0BWP7T $T=404720 137600 1 180 $X=402750 $Y=137365
X382 715 1 2 1377 INVD0BWP7T $T=420400 145440 0 180 $X=418430 $Y=141230
X383 713 1 2 716 INVD0BWP7T $T=420960 121920 0 180 $X=418990 $Y=117710
X384 708 1 2 1382 INVD0BWP7T $T=419840 153280 1 0 $X=419550 $Y=149070
X385 658 1 2 1380 INVD0BWP7T $T=422080 145440 0 180 $X=420110 $Y=141230
X386 1361 1 2 1379 INVD0BWP7T $T=422640 129760 0 180 $X=420670 $Y=125550
X387 723 1 2 724 INVD0BWP7T $T=423760 106240 0 0 $X=423470 $Y=106005
X388 721 1 2 1383 INVD0BWP7T $T=427120 153280 1 0 $X=426830 $Y=149070
X389 710 1 2 1386 INVD0BWP7T $T=443360 121920 0 180 $X=441390 $Y=117710
X390 171 105 1 2 BUFFD1P5BWP7T $T=90000 114080 1 180 $X=86910 $Y=113845
X391 1098 349 1 2 BUFFD1P5BWP7T $T=154400 153280 1 0 $X=154110 $Y=149070
X392 1178 1195 1 2 BUFFD1P5BWP7T $T=224400 137600 1 0 $X=224110 $Y=133390
X393 1327 630 1 2 BUFFD1P5BWP7T $T=366080 161120 0 180 $X=362990 $Y=156910
X394 764 766 1 2 BUFFD1P5BWP7T $T=445040 137600 0 0 $X=444750 $Y=137365
X395 786 530 1 2 BUFFD1P5BWP7T $T=466320 145440 0 180 $X=463230 $Y=141230
X396 1195 1 2 466 INVD3BWP7T $T=234480 137600 1 180 $X=230830 $Y=137365
X397 588 448 2 1 466 1291 593 MAOI22D0BWP7T $T=321280 114080 0 0 $X=320990 $Y=113845
X398 646 645 2 1 646 636 645 MAOI22D0BWP7T $T=367200 106240 1 180 $X=362990 $Y=106005
X399 704 1366 2 1 704 703 1366 MAOI22D0BWP7T $T=408080 161120 1 180 $X=403870 $Y=160885
X466 948 1 2 921 BUFFD1BWP7T $T=49120 145440 1 180 $X=46590 $Y=145205
X467 989 1 2 997 BUFFD1BWP7T $T=79920 121920 0 0 $X=79630 $Y=121685
X468 996 1 2 998 BUFFD1BWP7T $T=83840 137600 0 180 $X=81310 $Y=133390
X469 164 1 2 1000 BUFFD1BWP7T $T=82160 121920 0 0 $X=81870 $Y=121685
X470 1008 1 2 1012 BUFFD1BWP7T $T=93360 121920 1 0 $X=93070 $Y=117710
X471 1003 1 2 1013 BUFFD1BWP7T $T=93360 129760 1 0 $X=93070 $Y=125550
X472 1092 1 2 1100 BUFFD1BWP7T $T=142640 114080 0 0 $X=142350 $Y=113845
X473 324 1 2 1026 BUFFD1BWP7T $T=148800 129760 0 180 $X=146270 $Y=125550
X474 1116 1 2 1111 BUFFD1BWP7T $T=151600 137600 1 0 $X=151310 $Y=133390
X475 342 1 2 1110 BUFFD1BWP7T $T=154960 129760 1 180 $X=152430 $Y=129525
X476 370 1 2 1125 BUFFD1BWP7T $T=171760 114080 0 180 $X=169230 $Y=109870
X477 1127 1 2 1129 BUFFD1BWP7T $T=170080 121920 0 0 $X=169790 $Y=121685
X478 1124 1 2 1132 BUFFD1BWP7T $T=171200 129760 0 0 $X=170910 $Y=129525
X479 1153 1 2 1152 BUFFD1BWP7T $T=196400 114080 1 180 $X=193870 $Y=113845
X480 1155 1 2 1140 BUFFD1BWP7T $T=198080 114080 0 180 $X=195550 $Y=109870
X481 1179 1 2 1184 BUFFD1BWP7T $T=219920 153280 1 0 $X=219630 $Y=149070
X482 1255 1 2 1257 BUFFD1BWP7T $T=294400 137600 1 0 $X=294110 $Y=133390
X483 1274 1 2 567 BUFFD1BWP7T $T=306720 153280 1 0 $X=306430 $Y=149070
X484 574 1 2 577 BUFFD1BWP7T $T=310080 168960 1 0 $X=309790 $Y=164750
X485 1292 1 2 592 BUFFD1BWP7T $T=325200 121920 1 180 $X=322670 $Y=121685
X486 668 1 2 671 BUFFD1BWP7T $T=381200 168960 1 0 $X=380910 $Y=164750
X487 687 1 2 638 BUFFD1BWP7T $T=395200 121920 1 180 $X=392670 $Y=121685
X488 1358 1 2 1362 BUFFD1BWP7T $T=394080 145440 0 0 $X=393790 $Y=145205
X489 674 1 2 713 BUFFD1BWP7T $T=417040 153280 0 0 $X=416750 $Y=153045
X490 707 1 2 718 BUFFD1BWP7T $T=418720 106240 0 0 $X=418430 $Y=106005
X491 726 1 2 728 BUFFD1BWP7T $T=424880 114080 1 0 $X=424590 $Y=109870
X492 775 1 2 779 BUFFD1BWP7T $T=461280 145440 1 0 $X=460990 $Y=141230
X493 777 1 2 1388 BUFFD1BWP7T $T=461280 161120 0 0 $X=460990 $Y=160885
X494 776 1 2 778 BUFFD1BWP7T $T=461840 153280 1 0 $X=461550 $Y=149070
X495 1 2 DCAP4BWP7T $T=21120 114080 1 0 $X=20830 $Y=109870
X496 1 2 DCAP4BWP7T $T=21120 137600 1 0 $X=20830 $Y=133390
X497 1 2 DCAP4BWP7T $T=21120 153280 0 0 $X=20830 $Y=153045
X498 1 2 DCAP4BWP7T $T=42400 121920 0 0 $X=42110 $Y=121685
X499 1 2 DCAP4BWP7T $T=55280 145440 1 0 $X=54990 $Y=141230
X500 1 2 DCAP4BWP7T $T=64800 137600 1 0 $X=64510 $Y=133390
X501 1 2 DCAP4BWP7T $T=85520 145440 0 0 $X=85230 $Y=145205
X502 1 2 DCAP4BWP7T $T=86080 129760 0 0 $X=85790 $Y=129525
X503 1 2 DCAP4BWP7T $T=115760 153280 0 0 $X=115470 $Y=153045
X504 1 2 DCAP4BWP7T $T=152160 153280 1 0 $X=151870 $Y=149070
X505 1 2 DCAP4BWP7T $T=168400 161120 1 0 $X=168110 $Y=156910
X506 1 2 DCAP4BWP7T $T=170640 137600 1 0 $X=170350 $Y=133390
X507 1 2 DCAP4BWP7T $T=189680 129760 1 0 $X=189390 $Y=125550
X508 1 2 DCAP4BWP7T $T=199760 153280 0 0 $X=199470 $Y=153045
X509 1 2 DCAP4BWP7T $T=213760 145440 0 0 $X=213470 $Y=145205
X510 1 2 DCAP4BWP7T $T=217680 161120 0 0 $X=217390 $Y=160885
X511 1 2 DCAP4BWP7T $T=222160 137600 1 0 $X=221870 $Y=133390
X512 1 2 DCAP4BWP7T $T=222160 153280 1 0 $X=221870 $Y=149070
X513 1 2 DCAP4BWP7T $T=224960 153280 0 0 $X=224670 $Y=153045
X514 1 2 DCAP4BWP7T $T=231680 106240 0 0 $X=231390 $Y=106005
X515 1 2 DCAP4BWP7T $T=241760 121920 1 0 $X=241470 $Y=117710
X516 1 2 DCAP4BWP7T $T=260800 137600 1 0 $X=260510 $Y=133390
X517 1 2 DCAP4BWP7T $T=277600 106240 0 0 $X=277310 $Y=106005
X518 1 2 DCAP4BWP7T $T=303920 121920 1 0 $X=303630 $Y=117710
X519 1 2 DCAP4BWP7T $T=309520 129760 1 0 $X=309230 $Y=125550
X520 1 2 DCAP4BWP7T $T=325760 153280 1 0 $X=325470 $Y=149070
X521 1 2 DCAP4BWP7T $T=345360 129760 1 0 $X=345070 $Y=125550
X522 1 2 DCAP4BWP7T $T=345360 137600 1 0 $X=345070 $Y=133390
X523 1 2 DCAP4BWP7T $T=376720 106240 0 0 $X=376430 $Y=106005
X524 1 2 DCAP4BWP7T $T=378960 168960 1 0 $X=378670 $Y=164750
X525 1 2 DCAP4BWP7T $T=382320 121920 1 0 $X=382030 $Y=117710
X526 1 2 DCAP4BWP7T $T=389600 145440 0 0 $X=389310 $Y=145205
X527 1 2 DCAP4BWP7T $T=395200 161120 0 0 $X=394910 $Y=160885
X528 1 2 DCAP4BWP7T $T=396880 129760 0 0 $X=396590 $Y=129525
X529 1 2 DCAP4BWP7T $T=432720 145440 1 0 $X=432430 $Y=141230
X530 1 2 DCAP4BWP7T $T=471920 153280 0 0 $X=471630 $Y=153045
X531 1 2 ICV_3 $T=31200 114080 0 0 $X=30910 $Y=113845
X532 1 2 ICV_3 $T=31200 161120 1 0 $X=30910 $Y=156910
X533 1 2 ICV_3 $T=31200 168960 1 0 $X=30910 $Y=164750
X534 1 2 ICV_3 $T=35120 137600 0 0 $X=34830 $Y=137365
X535 1 2 ICV_3 $T=39600 129760 1 0 $X=39310 $Y=125550
X536 1 2 ICV_3 $T=39600 161120 1 0 $X=39310 $Y=156910
X537 1 2 ICV_3 $T=44080 145440 0 0 $X=43790 $Y=145205
X538 1 2 ICV_3 $T=62560 145440 0 0 $X=62270 $Y=145205
X539 1 2 ICV_3 $T=73200 106240 0 0 $X=72910 $Y=106005
X540 1 2 ICV_3 $T=73200 129760 1 0 $X=72910 $Y=125550
X541 1 2 ICV_3 $T=73200 129760 0 0 $X=72910 $Y=129525
X542 1 2 ICV_3 $T=77120 121920 0 0 $X=76830 $Y=121685
X543 1 2 ICV_3 $T=77120 153280 0 0 $X=76830 $Y=153045
X544 1 2 ICV_3 $T=77120 168960 1 0 $X=76830 $Y=164750
X545 1 2 ICV_3 $T=88880 168960 1 0 $X=88590 $Y=164750
X546 1 2 ICV_3 $T=94480 114080 1 0 $X=94190 $Y=109870
X547 1 2 ICV_3 $T=94480 121920 0 0 $X=94190 $Y=121685
X548 1 2 ICV_3 $T=103440 114080 1 0 $X=103150 $Y=109870
X549 1 2 ICV_3 $T=115200 137600 0 0 $X=114910 $Y=137365
X550 1 2 ICV_3 $T=115200 145440 1 0 $X=114910 $Y=141230
X551 1 2 ICV_3 $T=119120 114080 1 0 $X=118830 $Y=109870
X552 1 2 ICV_3 $T=119120 121920 1 0 $X=118830 $Y=117710
X553 1 2 ICV_3 $T=119120 121920 0 0 $X=118830 $Y=121685
X554 1 2 ICV_3 $T=119120 129760 1 0 $X=118830 $Y=125550
X555 1 2 ICV_3 $T=119120 161120 0 0 $X=118830 $Y=160885
X556 1 2 ICV_3 $T=125840 161120 0 0 $X=125550 $Y=160885
X557 1 2 ICV_3 $T=128080 161120 1 0 $X=127790 $Y=156910
X558 1 2 ICV_3 $T=135360 121920 0 0 $X=135070 $Y=121685
X559 1 2 ICV_3 $T=138720 129760 1 0 $X=138430 $Y=125550
X560 1 2 ICV_3 $T=147120 106240 0 0 $X=146830 $Y=106005
X561 1 2 ICV_3 $T=157200 121920 1 0 $X=156910 $Y=117710
X562 1 2 ICV_3 $T=157200 121920 0 0 $X=156910 $Y=121685
X563 1 2 ICV_3 $T=157200 137600 0 0 $X=156910 $Y=137365
X564 1 2 ICV_3 $T=157200 145440 0 0 $X=156910 $Y=145205
X565 1 2 ICV_3 $T=157200 153280 1 0 $X=156910 $Y=149070
X566 1 2 ICV_3 $T=157200 168960 1 0 $X=156910 $Y=164750
X567 1 2 ICV_3 $T=165600 129760 1 0 $X=165310 $Y=125550
X568 1 2 ICV_3 $T=165600 137600 0 0 $X=165310 $Y=137365
X569 1 2 ICV_3 $T=165600 153280 1 0 $X=165310 $Y=149070
X570 1 2 ICV_3 $T=186880 137600 0 0 $X=186590 $Y=137365
X571 1 2 ICV_3 $T=191360 121920 1 0 $X=191070 $Y=117710
X572 1 2 ICV_3 $T=199200 114080 0 0 $X=198910 $Y=113845
X573 1 2 ICV_3 $T=199200 137600 0 0 $X=198910 $Y=137365
X574 1 2 ICV_3 $T=199200 145440 1 0 $X=198910 $Y=141230
X575 1 2 ICV_3 $T=199200 161120 0 0 $X=198910 $Y=160885
X576 1 2 ICV_3 $T=207600 114080 1 0 $X=207310 $Y=109870
X577 1 2 ICV_3 $T=241200 114080 1 0 $X=240910 $Y=109870
X578 1 2 ICV_3 $T=241200 137600 1 0 $X=240910 $Y=133390
X579 1 2 ICV_3 $T=245120 145440 1 0 $X=244830 $Y=141230
X580 1 2 ICV_3 $T=249600 121920 1 0 $X=249310 $Y=117710
X581 1 2 ICV_3 $T=249600 129760 0 0 $X=249310 $Y=129525
X582 1 2 ICV_3 $T=249600 137600 0 0 $X=249310 $Y=137365
X583 1 2 ICV_3 $T=250720 161120 1 0 $X=250430 $Y=156910
X584 1 2 ICV_3 $T=258560 121920 1 0 $X=258270 $Y=117710
X585 1 2 ICV_3 $T=266960 145440 1 0 $X=266670 $Y=141230
X586 1 2 ICV_3 $T=269760 145440 0 0 $X=269470 $Y=145205
X587 1 2 ICV_3 $T=273120 121920 1 0 $X=272830 $Y=117710
X588 1 2 ICV_3 $T=283200 137600 1 0 $X=282910 $Y=133390
X589 1 2 ICV_3 $T=283200 153280 0 0 $X=282910 $Y=153045
X590 1 2 ICV_3 $T=287120 161120 0 0 $X=286830 $Y=160885
X591 1 2 ICV_3 $T=291600 137600 1 0 $X=291310 $Y=133390
X592 1 2 ICV_3 $T=303920 153280 1 0 $X=303630 $Y=149070
X593 1 2 ICV_3 $T=314560 114080 1 0 $X=314270 $Y=109870
X594 1 2 ICV_3 $T=325200 114080 0 0 $X=324910 $Y=113845
X595 1 2 ICV_3 $T=325200 121920 0 0 $X=324910 $Y=121685
X596 1 2 ICV_3 $T=325200 137600 1 0 $X=324910 $Y=133390
X597 1 2 ICV_3 $T=325200 161120 1 0 $X=324910 $Y=156910
X598 1 2 ICV_3 $T=325200 168960 1 0 $X=324910 $Y=164750
X599 1 2 ICV_3 $T=343680 161120 1 0 $X=343390 $Y=156910
X600 1 2 ICV_3 $T=352640 114080 1 0 $X=352350 $Y=109870
X601 1 2 ICV_3 $T=354880 168960 1 0 $X=354590 $Y=164750
X602 1 2 ICV_3 $T=367200 106240 0 0 $X=366910 $Y=106005
X603 1 2 ICV_3 $T=367200 114080 0 0 $X=366910 $Y=113845
X604 1 2 ICV_3 $T=367200 121920 1 0 $X=366910 $Y=117710
X605 1 2 ICV_3 $T=386800 129760 1 0 $X=386510 $Y=125550
X606 1 2 ICV_3 $T=390720 114080 0 0 $X=390430 $Y=113845
X607 1 2 ICV_3 $T=403600 145440 0 0 $X=403310 $Y=145205
X608 1 2 ICV_3 $T=409200 106240 0 0 $X=408910 $Y=106005
X609 1 2 ICV_3 $T=409200 121920 0 0 $X=408910 $Y=121685
X610 1 2 ICV_3 $T=420960 106240 0 0 $X=420670 $Y=106005
X611 1 2 ICV_3 $T=422080 114080 1 0 $X=421790 $Y=109870
X612 1 2 ICV_3 $T=438880 121920 1 0 $X=438590 $Y=117710
X613 1 2 ICV_3 $T=451200 145440 0 0 $X=450910 $Y=145205
X614 1 2 ICV_3 $T=471360 121920 1 0 $X=471070 $Y=117710
X615 1 2 ICV_3 $T=471360 137600 1 0 $X=471070 $Y=133390
X616 1 2 ICV_3 $T=471360 153280 1 0 $X=471070 $Y=149070
X617 1 2 DCAP8BWP7T $T=26720 161120 1 0 $X=26430 $Y=156910
X618 1 2 DCAP8BWP7T $T=26720 168960 1 0 $X=26430 $Y=164750
X619 1 2 DCAP8BWP7T $T=27840 161120 0 0 $X=27550 $Y=160885
X620 1 2 DCAP8BWP7T $T=35120 137600 1 0 $X=34830 $Y=133390
X621 1 2 DCAP8BWP7T $T=58080 145440 0 0 $X=57790 $Y=145205
X622 1 2 DCAP8BWP7T $T=62000 114080 1 0 $X=61710 $Y=109870
X623 1 2 DCAP8BWP7T $T=63120 161120 0 0 $X=62830 $Y=160885
X624 1 2 DCAP8BWP7T $T=77120 153280 1 0 $X=76830 $Y=149070
X625 1 2 DCAP8BWP7T $T=90560 129760 0 0 $X=90270 $Y=129525
X626 1 2 DCAP8BWP7T $T=91680 145440 0 0 $X=91390 $Y=145205
X627 1 2 DCAP8BWP7T $T=98960 153280 1 0 $X=98670 $Y=149070
X628 1 2 DCAP8BWP7T $T=110720 137600 0 0 $X=110430 $Y=137365
X629 1 2 DCAP8BWP7T $T=111840 114080 0 0 $X=111550 $Y=113845
X630 1 2 DCAP8BWP7T $T=111840 129760 1 0 $X=111550 $Y=125550
X631 1 2 DCAP8BWP7T $T=123600 145440 1 0 $X=123310 $Y=141230
X632 1 2 DCAP8BWP7T $T=124160 121920 1 0 $X=123870 $Y=117710
X633 1 2 DCAP8BWP7T $T=129200 145440 0 0 $X=128910 $Y=145205
X634 1 2 DCAP8BWP7T $T=135920 137600 1 0 $X=135630 $Y=133390
X635 1 2 DCAP8BWP7T $T=142640 161120 0 0 $X=142350 $Y=160885
X636 1 2 DCAP8BWP7T $T=145440 153280 0 0 $X=145150 $Y=153045
X637 1 2 DCAP8BWP7T $T=146560 129760 0 0 $X=146270 $Y=129525
X638 1 2 DCAP8BWP7T $T=147120 168960 1 0 $X=146830 $Y=164750
X639 1 2 DCAP8BWP7T $T=153840 137600 1 0 $X=153550 $Y=133390
X640 1 2 DCAP8BWP7T $T=155520 114080 1 0 $X=155230 $Y=109870
X641 1 2 DCAP8BWP7T $T=161120 153280 0 0 $X=160830 $Y=153045
X642 1 2 DCAP8BWP7T $T=173440 129760 0 0 $X=173150 $Y=129525
X643 1 2 DCAP8BWP7T $T=177360 153280 0 0 $X=177070 $Y=153045
X644 1 2 DCAP8BWP7T $T=182400 129760 0 0 $X=182110 $Y=129525
X645 1 2 DCAP8BWP7T $T=189680 114080 0 0 $X=189390 $Y=113845
X646 1 2 DCAP8BWP7T $T=194160 129760 1 0 $X=193870 $Y=125550
X647 1 2 DCAP8BWP7T $T=194160 137600 1 0 $X=193870 $Y=133390
X648 1 2 DCAP8BWP7T $T=194720 137600 0 0 $X=194430 $Y=137365
X649 1 2 DCAP8BWP7T $T=194720 161120 0 0 $X=194430 $Y=160885
X650 1 2 DCAP8BWP7T $T=209840 153280 1 0 $X=209550 $Y=149070
X651 1 2 DCAP8BWP7T $T=211520 145440 1 0 $X=211230 $Y=141230
X652 1 2 DCAP8BWP7T $T=213200 121920 1 0 $X=212910 $Y=117710
X653 1 2 DCAP8BWP7T $T=226640 153280 1 0 $X=226350 $Y=149070
X654 1 2 DCAP8BWP7T $T=230560 153280 0 0 $X=230270 $Y=153045
X655 1 2 DCAP8BWP7T $T=236160 129760 0 0 $X=235870 $Y=129525
X656 1 2 DCAP8BWP7T $T=236720 114080 1 0 $X=236430 $Y=109870
X657 1 2 DCAP8BWP7T $T=237840 145440 1 0 $X=237550 $Y=141230
X658 1 2 DCAP8BWP7T $T=237840 153280 1 0 $X=237550 $Y=149070
X659 1 2 DCAP8BWP7T $T=238960 145440 0 0 $X=238670 $Y=145205
X660 1 2 DCAP8BWP7T $T=239520 106240 0 0 $X=239230 $Y=106005
X661 1 2 DCAP8BWP7T $T=245120 137600 0 0 $X=244830 $Y=137365
X662 1 2 DCAP8BWP7T $T=251280 114080 0 0 $X=250990 $Y=113845
X663 1 2 DCAP8BWP7T $T=264720 161120 0 0 $X=264430 $Y=160885
X664 1 2 DCAP8BWP7T $T=265280 153280 1 0 $X=264990 $Y=149070
X665 1 2 DCAP8BWP7T $T=270880 106240 0 0 $X=270590 $Y=106005
X666 1 2 DCAP8BWP7T $T=279840 121920 0 0 $X=279550 $Y=121685
X667 1 2 DCAP8BWP7T $T=279840 161120 0 0 $X=279550 $Y=160885
X668 1 2 DCAP8BWP7T $T=281520 145440 0 0 $X=281230 $Y=145205
X669 1 2 DCAP8BWP7T $T=287120 129760 1 0 $X=286830 $Y=125550
X670 1 2 DCAP8BWP7T $T=294400 153280 0 0 $X=294110 $Y=153045
X671 1 2 DCAP8BWP7T $T=297760 129760 1 0 $X=297470 $Y=125550
X672 1 2 DCAP8BWP7T $T=299440 137600 1 0 $X=299150 $Y=133390
X673 1 2 DCAP8BWP7T $T=300560 137600 0 0 $X=300270 $Y=137365
X674 1 2 DCAP8BWP7T $T=302800 161120 1 0 $X=302510 $Y=156910
X675 1 2 DCAP8BWP7T $T=308400 137600 0 0 $X=308110 $Y=137365
X676 1 2 DCAP8BWP7T $T=312320 161120 0 0 $X=312030 $Y=160885
X677 1 2 DCAP8BWP7T $T=319040 161120 1 0 $X=318750 $Y=156910
X678 1 2 DCAP8BWP7T $T=322960 145440 1 0 $X=322670 $Y=141230
X679 1 2 DCAP8BWP7T $T=323520 106240 0 0 $X=323230 $Y=106005
X680 1 2 DCAP8BWP7T $T=336400 114080 0 0 $X=336110 $Y=113845
X681 1 2 DCAP8BWP7T $T=340320 153280 0 0 $X=340030 $Y=153045
X682 1 2 DCAP8BWP7T $T=347040 114080 0 0 $X=346750 $Y=113845
X683 1 2 DCAP8BWP7T $T=350400 168960 1 0 $X=350110 $Y=164750
X684 1 2 DCAP8BWP7T $T=362160 137600 0 0 $X=361870 $Y=137365
X685 1 2 DCAP8BWP7T $T=362160 153280 0 0 $X=361870 $Y=153045
X686 1 2 DCAP8BWP7T $T=364960 129760 0 0 $X=364670 $Y=129525
X687 1 2 DCAP8BWP7T $T=371120 168960 1 0 $X=370830 $Y=164750
X688 1 2 DCAP8BWP7T $T=376720 137600 1 0 $X=376430 $Y=133390
X689 1 2 DCAP8BWP7T $T=384560 137600 1 0 $X=384270 $Y=133390
X690 1 2 DCAP8BWP7T $T=384560 145440 1 0 $X=384270 $Y=141230
X691 1 2 DCAP8BWP7T $T=386240 114080 0 0 $X=385950 $Y=113845
X692 1 2 DCAP8BWP7T $T=390160 121920 1 0 $X=389870 $Y=117710
X693 1 2 DCAP8BWP7T $T=395200 121920 0 0 $X=394910 $Y=121685
X694 1 2 DCAP8BWP7T $T=399120 161120 0 0 $X=398830 $Y=160885
X695 1 2 DCAP8BWP7T $T=404160 129760 1 0 $X=403870 $Y=125550
X696 1 2 DCAP8BWP7T $T=404160 153280 0 0 $X=403870 $Y=153045
X697 1 2 DCAP8BWP7T $T=404720 106240 0 0 $X=404430 $Y=106005
X698 1 2 DCAP8BWP7T $T=404720 121920 0 0 $X=404430 $Y=121685
X699 1 2 DCAP8BWP7T $T=404720 137600 0 0 $X=404430 $Y=137365
X700 1 2 DCAP8BWP7T $T=407520 121920 1 0 $X=407230 $Y=117710
X701 1 2 DCAP8BWP7T $T=423200 137600 0 0 $X=422910 $Y=137365
X702 1 2 DCAP8BWP7T $T=425440 106240 0 0 $X=425150 $Y=106005
X703 1 2 DCAP8BWP7T $T=426560 129760 0 0 $X=426270 $Y=129525
X704 1 2 DCAP8BWP7T $T=431040 137600 1 0 $X=430750 $Y=133390
X705 1 2 DCAP8BWP7T $T=432160 168960 1 0 $X=431870 $Y=164750
X706 1 2 DCAP8BWP7T $T=437760 137600 1 0 $X=437470 $Y=133390
X707 1 2 DCAP8BWP7T $T=440560 137600 0 0 $X=440270 $Y=137365
X708 1 2 DCAP8BWP7T $T=446160 106240 0 0 $X=445870 $Y=106005
X709 1 2 DCAP8BWP7T $T=446720 145440 0 0 $X=446430 $Y=145205
X710 1 2 DCAP8BWP7T $T=447840 137600 1 0 $X=447550 $Y=133390
X711 1 2 DCAP8BWP7T $T=447840 137600 0 0 $X=447550 $Y=137365
X712 1 2 DCAP8BWP7T $T=447840 161120 0 0 $X=447550 $Y=160885
X713 1 2 DCAP8BWP7T $T=466320 145440 1 0 $X=466030 $Y=141230
X714 1 2 DCAP8BWP7T $T=466880 153280 1 0 $X=466590 $Y=149070
X715 2 1 DCAPBWP7T $T=25040 137600 1 0 $X=24750 $Y=133390
X716 2 1 DCAPBWP7T $T=67600 161120 0 0 $X=67310 $Y=160885
X717 2 1 DCAPBWP7T $T=69840 129760 1 0 $X=69550 $Y=125550
X718 2 1 DCAPBWP7T $T=81600 153280 1 0 $X=81310 $Y=149070
X719 2 1 DCAPBWP7T $T=90560 114080 1 0 $X=90270 $Y=109870
X720 2 1 DCAPBWP7T $T=93920 137600 0 0 $X=93630 $Y=137365
X721 2 1 DCAPBWP7T $T=96160 145440 0 0 $X=95870 $Y=145205
X722 2 1 DCAPBWP7T $T=105680 137600 0 0 $X=105390 $Y=137365
X723 2 1 DCAPBWP7T $T=111840 161120 0 0 $X=111550 $Y=160885
X724 2 1 DCAPBWP7T $T=126960 153280 1 0 $X=126670 $Y=149070
X725 2 1 DCAPBWP7T $T=128080 145440 1 0 $X=127790 $Y=141230
X726 2 1 DCAPBWP7T $T=151040 129760 0 0 $X=150750 $Y=129525
X727 2 1 DCAPBWP7T $T=165600 153280 0 0 $X=165310 $Y=153045
X728 2 1 DCAPBWP7T $T=171200 153280 0 0 $X=170910 $Y=153045
X729 2 1 DCAPBWP7T $T=174560 168960 1 0 $X=174270 $Y=164750
X730 2 1 DCAPBWP7T $T=176240 145440 1 0 $X=175950 $Y=141230
X731 2 1 DCAPBWP7T $T=182400 114080 1 0 $X=182110 $Y=109870
X732 2 1 DCAPBWP7T $T=200320 121920 0 0 $X=200030 $Y=121685
X733 2 1 DCAPBWP7T $T=200320 145440 0 0 $X=200030 $Y=145205
X734 2 1 DCAPBWP7T $T=232800 145440 1 0 $X=232510 $Y=141230
X735 2 1 DCAPBWP7T $T=242320 129760 1 0 $X=242030 $Y=125550
X736 2 1 DCAPBWP7T $T=249600 106240 0 0 $X=249310 $Y=106005
X737 2 1 DCAPBWP7T $T=249600 114080 1 0 $X=249310 $Y=109870
X738 2 1 DCAPBWP7T $T=261920 114080 0 0 $X=261630 $Y=113845
X739 2 1 DCAPBWP7T $T=269760 129760 0 0 $X=269470 $Y=129525
X740 2 1 DCAPBWP7T $T=270320 153280 0 0 $X=270030 $Y=153045
X741 2 1 DCAPBWP7T $T=296080 161120 1 0 $X=295790 $Y=156910
X742 2 1 DCAPBWP7T $T=305040 137600 0 0 $X=304750 $Y=137365
X743 2 1 DCAPBWP7T $T=307280 114080 1 0 $X=306990 $Y=109870
X744 2 1 DCAPBWP7T $T=317920 137600 0 0 $X=317630 $Y=137365
X745 2 1 DCAPBWP7T $T=333600 121920 1 0 $X=333310 $Y=117710
X746 2 1 DCAPBWP7T $T=333600 129760 1 0 $X=333310 $Y=125550
X747 2 1 DCAPBWP7T $T=333600 161120 1 0 $X=333310 $Y=156910
X748 2 1 DCAPBWP7T $T=342000 114080 1 0 $X=341710 $Y=109870
X749 2 1 DCAPBWP7T $T=377840 114080 1 0 $X=377550 $Y=109870
X750 2 1 DCAPBWP7T $T=384560 153280 1 0 $X=384270 $Y=149070
X751 2 1 DCAPBWP7T $T=389040 137600 1 0 $X=388750 $Y=133390
X752 2 1 DCAPBWP7T $T=394640 121920 1 0 $X=394350 $Y=117710
X753 2 1 DCAPBWP7T $T=399680 121920 0 0 $X=399390 $Y=121685
X754 2 1 DCAPBWP7T $T=410320 137600 1 0 $X=410030 $Y=133390
X755 2 1 DCAPBWP7T $T=431040 129760 0 0 $X=430750 $Y=129525
X756 2 1 DCAPBWP7T $T=436640 168960 1 0 $X=436350 $Y=164750
X757 2 1 DCAPBWP7T $T=452320 114080 1 0 $X=452030 $Y=109870
X758 2 1 DCAPBWP7T $T=452320 129760 1 0 $X=452030 $Y=125550
X759 2 1 DCAPBWP7T $T=452320 137600 0 0 $X=452030 $Y=137365
X760 2 1 DCAPBWP7T $T=452320 145440 1 0 $X=452030 $Y=141230
X761 2 1 DCAPBWP7T $T=459600 129760 0 0 $X=459310 $Y=129525
X762 2 1 DCAPBWP7T $T=459600 145440 1 0 $X=459310 $Y=141230
X763 627 625 608 572 1295 613 1 2 617 AO222D1BWP7T $T=350400 168960 0 180 $X=343390 $Y=164750
X764 1 2 ICV_4 $T=30080 129760 0 0 $X=29790 $Y=129525
X765 1 2 ICV_4 $T=55280 168960 1 0 $X=54990 $Y=164750
X766 1 2 ICV_4 $T=72080 137600 0 0 $X=71790 $Y=137365
X767 1 2 ICV_4 $T=119120 137600 0 0 $X=118830 $Y=137365
X768 1 2 ICV_4 $T=119120 168960 1 0 $X=118830 $Y=164750
X769 1 2 ICV_4 $T=156080 129760 1 0 $X=155790 $Y=125550
X770 1 2 ICV_4 $T=156080 161120 1 0 $X=155790 $Y=156910
X771 1 2 ICV_4 $T=161120 168960 1 0 $X=160830 $Y=164750
X772 1 2 ICV_4 $T=185760 153280 0 0 $X=185470 $Y=153045
X773 1 2 ICV_4 $T=186880 153280 1 0 $X=186590 $Y=149070
X774 1 2 ICV_4 $T=198080 114080 1 0 $X=197790 $Y=109870
X775 1 2 ICV_4 $T=203120 145440 1 0 $X=202830 $Y=141230
X776 1 2 ICV_4 $T=245120 114080 0 0 $X=244830 $Y=113845
X777 1 2 ICV_4 $T=245120 121920 0 0 $X=244830 $Y=121685
X778 1 2 ICV_4 $T=255760 168960 1 0 $X=255470 $Y=164750
X779 1 2 ICV_4 $T=265840 114080 1 0 $X=265550 $Y=109870
X780 1 2 ICV_4 $T=272560 168960 1 0 $X=272270 $Y=164750
X781 1 2 ICV_4 $T=273680 129760 1 0 $X=273390 $Y=125550
X782 1 2 ICV_4 $T=282080 137600 0 0 $X=281790 $Y=137365
X783 1 2 ICV_4 $T=282080 161120 1 0 $X=281790 $Y=156910
X784 1 2 ICV_4 $T=287120 121920 0 0 $X=286830 $Y=121685
X785 1 2 ICV_4 $T=293840 106240 0 0 $X=293550 $Y=106005
X786 1 2 ICV_4 $T=296080 153280 1 0 $X=295790 $Y=149070
X787 1 2 ICV_4 $T=324080 121920 1 0 $X=323790 $Y=117710
X788 1 2 ICV_4 $T=338080 153280 1 0 $X=337790 $Y=149070
X789 1 2 ICV_4 $T=339760 121920 1 0 $X=339470 $Y=117710
X790 1 2 ICV_4 $T=339760 137600 1 0 $X=339470 $Y=133390
X791 1 2 ICV_4 $T=366080 137600 1 0 $X=365790 $Y=133390
X792 1 2 ICV_4 $T=366080 161120 1 0 $X=365790 $Y=156910
X793 1 2 ICV_4 $T=387360 168960 1 0 $X=387070 $Y=164750
X794 1 2 ICV_4 $T=399120 106240 0 0 $X=398830 $Y=106005
X795 1 2 ICV_4 $T=408080 129760 0 0 $X=407790 $Y=129525
X796 1 2 ICV_4 $T=408080 145440 0 0 $X=407790 $Y=145205
X797 1 2 ICV_4 $T=408080 153280 1 0 $X=407790 $Y=149070
X798 1 2 ICV_4 $T=413120 114080 0 0 $X=412830 $Y=113845
X799 1 2 ICV_4 $T=413120 153280 0 0 $X=412830 $Y=153045
X800 1 2 ICV_4 $T=450080 129760 0 0 $X=449790 $Y=129525
X801 1 2 ICV_4 $T=455120 153280 0 0 $X=454830 $Y=153045
X802 374 677 525 2 1 624 DFCNQD1BWP7T $T=392960 121920 1 180 $X=380350 $Y=121685
X803 374 725 525 2 1 707 DFCNQD1BWP7T $T=428240 121920 1 180 $X=415630 $Y=121685
X1067 1 2 ICV_8 $T=20000 129760 1 0 $X=19710 $Y=125550
X1068 1 2 ICV_8 $T=20000 153280 1 0 $X=19710 $Y=149070
X1069 1 2 ICV_8 $T=20000 161120 0 0 $X=19710 $Y=160885
X1070 1 2 ICV_8 $T=34000 114080 0 0 $X=33710 $Y=113845
X1071 1 2 ICV_8 $T=34000 121920 1 0 $X=33710 $Y=117710
X1072 1 2 ICV_8 $T=34000 129760 0 0 $X=33710 $Y=129525
X1073 1 2 ICV_8 $T=34000 145440 0 0 $X=33710 $Y=145205
X1074 1 2 ICV_8 $T=76000 129760 1 0 $X=75710 $Y=125550
X1075 1 2 ICV_8 $T=76000 145440 0 0 $X=75710 $Y=145205
X1076 1 2 ICV_8 $T=118000 106240 0 0 $X=117710 $Y=106005
X1077 1 2 ICV_8 $T=118000 137600 1 0 $X=117710 $Y=133390
X1078 1 2 ICV_8 $T=118000 145440 1 0 $X=117710 $Y=141230
X1079 1 2 ICV_8 $T=118000 153280 0 0 $X=117710 $Y=153045
X1080 1 2 ICV_8 $T=160000 161120 1 0 $X=159710 $Y=156910
X1081 1 2 ICV_8 $T=202000 114080 0 0 $X=201710 $Y=113845
X1082 1 2 ICV_8 $T=202000 153280 1 0 $X=201710 $Y=149070
X1083 1 2 ICV_8 $T=202000 168960 1 0 $X=201710 $Y=164750
X1084 1 2 ICV_8 $T=244000 137600 1 0 $X=243710 $Y=133390
X1085 1 2 ICV_8 $T=286000 145440 1 0 $X=285710 $Y=141230
X1086 1 2 ICV_8 $T=286000 145440 0 0 $X=285710 $Y=145205
X1087 1 2 ICV_8 $T=328000 106240 0 0 $X=327710 $Y=106005
X1088 1 2 ICV_8 $T=328000 137600 1 0 $X=327710 $Y=133390
X1089 1 2 ICV_8 $T=328000 153280 0 0 $X=327710 $Y=153045
X1090 1 2 ICV_8 $T=370000 106240 0 0 $X=369710 $Y=106005
X1091 1 2 ICV_8 $T=370000 161120 0 0 $X=369710 $Y=160885
X1092 1 2 ICV_8 $T=412000 121920 0 0 $X=411710 $Y=121685
X1093 1 2 ICV_8 $T=454000 145440 0 0 $X=453710 $Y=145205
X1094 1 2 ICV_9 $T=34000 129760 1 0 $X=33710 $Y=125550
X1095 1 2 ICV_9 $T=34000 161120 1 0 $X=33710 $Y=156910
X1096 1 2 ICV_9 $T=34000 168960 1 0 $X=33710 $Y=164750
X1097 1 2 ICV_9 $T=76000 106240 0 0 $X=75710 $Y=106005
X1098 1 2 ICV_9 $T=76000 137600 1 0 $X=75710 $Y=133390
X1099 1 2 ICV_9 $T=76000 145440 1 0 $X=75710 $Y=141230
X1100 1 2 ICV_9 $T=76000 161120 1 0 $X=75710 $Y=156910
X1101 1 2 ICV_9 $T=118000 161120 1 0 $X=117710 $Y=156910
X1102 1 2 ICV_9 $T=160000 114080 1 0 $X=159710 $Y=109870
X1103 1 2 ICV_9 $T=160000 129760 1 0 $X=159710 $Y=125550
X1104 1 2 ICV_9 $T=160000 137600 0 0 $X=159710 $Y=137365
X1105 1 2 ICV_9 $T=160000 145440 1 0 $X=159710 $Y=141230
X1106 1 2 ICV_9 $T=160000 145440 0 0 $X=159710 $Y=145205
X1107 1 2 ICV_9 $T=160000 153280 1 0 $X=159710 $Y=149070
X1108 1 2 ICV_9 $T=160000 161120 0 0 $X=159710 $Y=160885
X1109 1 2 ICV_9 $T=202000 114080 1 0 $X=201710 $Y=109870
X1110 1 2 ICV_9 $T=202000 121920 1 0 $X=201710 $Y=117710
X1111 1 2 ICV_9 $T=202000 121920 0 0 $X=201710 $Y=121685
X1112 1 2 ICV_9 $T=202000 137600 1 0 $X=201710 $Y=133390
X1113 1 2 ICV_9 $T=202000 137600 0 0 $X=201710 $Y=137365
X1114 1 2 ICV_9 $T=202000 145440 0 0 $X=201710 $Y=145205
X1115 1 2 ICV_9 $T=244000 106240 0 0 $X=243710 $Y=106005
X1116 1 2 ICV_9 $T=244000 114080 1 0 $X=243710 $Y=109870
X1117 1 2 ICV_9 $T=244000 121920 1 0 $X=243710 $Y=117710
X1118 1 2 ICV_9 $T=244000 129760 1 0 $X=243710 $Y=125550
X1119 1 2 ICV_9 $T=244000 129760 0 0 $X=243710 $Y=129525
X1120 1 2 ICV_9 $T=244000 153280 0 0 $X=243710 $Y=153045
X1121 1 2 ICV_9 $T=244000 161120 0 0 $X=243710 $Y=160885
X1122 1 2 ICV_9 $T=286000 114080 1 0 $X=285710 $Y=109870
X1123 1 2 ICV_9 $T=286000 137600 1 0 $X=285710 $Y=133390
X1124 1 2 ICV_9 $T=286000 153280 1 0 $X=285710 $Y=149070
X1125 1 2 ICV_9 $T=328000 114080 1 0 $X=327710 $Y=109870
X1126 1 2 ICV_9 $T=328000 121920 1 0 $X=327710 $Y=117710
X1127 1 2 ICV_9 $T=328000 129760 1 0 $X=327710 $Y=125550
X1128 1 2 ICV_9 $T=328000 161120 1 0 $X=327710 $Y=156910
X1129 1 2 ICV_9 $T=328000 161120 0 0 $X=327710 $Y=160885
X1130 1 2 ICV_9 $T=328000 168960 1 0 $X=327710 $Y=164750
X1131 1 2 ICV_9 $T=370000 145440 1 0 $X=369710 $Y=141230
X1132 1 2 ICV_9 $T=370000 161120 1 0 $X=369710 $Y=156910
X1133 1 2 ICV_9 $T=412000 106240 0 0 $X=411710 $Y=106005
X1134 1 2 ICV_9 $T=412000 114080 1 0 $X=411710 $Y=109870
X1135 1 2 ICV_9 $T=412000 129760 1 0 $X=411710 $Y=125550
X1136 1 2 ICV_9 $T=412000 137600 1 0 $X=411710 $Y=133390
X1137 1 2 ICV_9 $T=412000 168960 1 0 $X=411710 $Y=164750
X1138 1 2 ICV_9 $T=454000 114080 1 0 $X=453710 $Y=109870
X1139 1 2 ICV_9 $T=454000 129760 1 0 $X=453710 $Y=125550
X1140 1 2 ICV_9 $T=454000 129760 0 0 $X=453710 $Y=129525
X1141 1 2 ICV_9 $T=454000 137600 0 0 $X=453710 $Y=137365
X1142 1 2 ICV_9 $T=454000 145440 1 0 $X=453710 $Y=141230
X1182 1 2 ICV_13 $T=21120 114080 0 0 $X=20830 $Y=113845
X1183 1 2 ICV_13 $T=21120 161120 1 0 $X=20830 $Y=156910
X1184 1 2 ICV_13 $T=30640 129760 1 0 $X=30350 $Y=125550
X1185 1 2 ICV_13 $T=30640 145440 0 0 $X=30350 $Y=145205
X1186 1 2 ICV_13 $T=35120 121920 0 0 $X=34830 $Y=121685
X1187 1 2 ICV_13 $T=35120 145440 1 0 $X=34830 $Y=141230
X1188 1 2 ICV_13 $T=35120 153280 0 0 $X=34830 $Y=153045
X1189 1 2 ICV_13 $T=59200 137600 0 0 $X=58910 $Y=137365
X1190 1 2 ICV_13 $T=60880 121920 1 0 $X=60590 $Y=117710
X1191 1 2 ICV_13 $T=64240 168960 1 0 $X=63950 $Y=164750
X1192 1 2 ICV_13 $T=66480 114080 1 0 $X=66190 $Y=109870
X1193 1 2 ICV_13 $T=66480 137600 0 0 $X=66190 $Y=137365
X1194 1 2 ICV_13 $T=77120 114080 0 0 $X=76830 $Y=113845
X1195 1 2 ICV_13 $T=77120 137600 0 0 $X=76830 $Y=137365
X1196 1 2 ICV_13 $T=81600 106240 0 0 $X=81310 $Y=106005
X1197 1 2 ICV_13 $T=98960 137600 0 0 $X=98670 $Y=137365
X1198 1 2 ICV_13 $T=100080 137600 1 0 $X=99790 $Y=133390
X1199 1 2 ICV_13 $T=103440 153280 1 0 $X=103150 $Y=149070
X1200 1 2 ICV_13 $T=114640 137600 1 0 $X=114350 $Y=133390
X1201 1 2 ICV_13 $T=114640 153280 1 0 $X=114350 $Y=149070
X1202 1 2 ICV_13 $T=114640 161120 1 0 $X=114350 $Y=156910
X1203 1 2 ICV_13 $T=119120 153280 1 0 $X=118830 $Y=149070
X1204 1 2 ICV_13 $T=126960 168960 1 0 $X=126670 $Y=164750
X1205 1 2 ICV_13 $T=131440 153280 0 0 $X=131150 $Y=153045
X1206 1 2 ICV_13 $T=133120 129760 0 0 $X=132830 $Y=129525
X1207 1 2 ICV_13 $T=138720 153280 0 0 $X=138430 $Y=153045
X1208 1 2 ICV_13 $T=156640 129760 0 0 $X=156350 $Y=129525
X1209 1 2 ICV_13 $T=156640 145440 1 0 $X=156350 $Y=141230
X1210 1 2 ICV_13 $T=156640 161120 0 0 $X=156350 $Y=160885
X1211 1 2 ICV_13 $T=161120 106240 0 0 $X=160830 $Y=106005
X1212 1 2 ICV_13 $T=161120 121920 1 0 $X=160830 $Y=117710
X1213 1 2 ICV_13 $T=161120 137600 1 0 $X=160830 $Y=133390
X1214 1 2 ICV_13 $T=165600 114080 1 0 $X=165310 $Y=109870
X1215 1 2 ICV_13 $T=171760 114080 1 0 $X=171470 $Y=109870
X1216 1 2 ICV_13 $T=172320 145440 0 0 $X=172030 $Y=145205
X1217 1 2 ICV_13 $T=175680 106240 0 0 $X=175390 $Y=106005
X1218 1 2 ICV_13 $T=180720 145440 0 0 $X=180430 $Y=145205
X1219 1 2 ICV_13 $T=187440 114080 1 0 $X=187150 $Y=109870
X1220 1 2 ICV_13 $T=198640 129760 1 0 $X=198350 $Y=125550
X1221 1 2 ICV_13 $T=198640 137600 1 0 $X=198350 $Y=133390
X1222 1 2 ICV_13 $T=198640 153280 1 0 $X=198350 $Y=149070
X1223 1 2 ICV_13 $T=203120 161120 0 0 $X=202830 $Y=160885
X1224 1 2 ICV_13 $T=207600 137600 0 0 $X=207310 $Y=137365
X1225 1 2 ICV_13 $T=227200 137600 0 0 $X=226910 $Y=137365
X1226 1 2 ICV_13 $T=240640 129760 0 0 $X=240350 $Y=129525
X1227 1 2 ICV_13 $T=245120 145440 0 0 $X=244830 $Y=145205
X1228 1 2 ICV_13 $T=245120 161120 1 0 $X=244830 $Y=156910
X1229 1 2 ICV_13 $T=245120 168960 1 0 $X=244830 $Y=164750
X1230 1 2 ICV_13 $T=249600 129760 1 0 $X=249310 $Y=125550
X1231 1 2 ICV_13 $T=255760 145440 0 0 $X=255470 $Y=145205
X1232 1 2 ICV_13 $T=282640 106240 0 0 $X=282350 $Y=106005
X1233 1 2 ICV_13 $T=282640 145440 1 0 $X=282350 $Y=141230
X1234 1 2 ICV_13 $T=287120 106240 0 0 $X=286830 $Y=106005
X1235 1 2 ICV_13 $T=287120 137600 0 0 $X=286830 $Y=137365
X1236 1 2 ICV_13 $T=287120 153280 0 0 $X=286830 $Y=153045
X1237 1 2 ICV_13 $T=291600 129760 1 0 $X=291310 $Y=125550
X1238 1 2 ICV_13 $T=302240 153280 0 0 $X=301950 $Y=153045
X1239 1 2 ICV_13 $T=312880 129760 0 0 $X=312590 $Y=129525
X1240 1 2 ICV_13 $T=316800 137600 1 0 $X=316510 $Y=133390
X1241 1 2 ICV_13 $T=324640 129760 1 0 $X=324350 $Y=125550
X1242 1 2 ICV_13 $T=324640 137600 0 0 $X=324350 $Y=137365
X1243 1 2 ICV_13 $T=329120 114080 0 0 $X=328830 $Y=113845
X1244 1 2 ICV_13 $T=329120 137600 0 0 $X=328830 $Y=137365
X1245 1 2 ICV_13 $T=333600 161120 0 0 $X=333310 $Y=160885
X1246 1 2 ICV_13 $T=338080 106240 0 0 $X=337790 $Y=106005
X1247 1 2 ICV_13 $T=338080 161120 1 0 $X=337790 $Y=156910
X1248 1 2 ICV_13 $T=340880 114080 0 0 $X=340590 $Y=113845
X1249 1 2 ICV_13 $T=356000 114080 0 0 $X=355710 $Y=113845
X1250 1 2 ICV_13 $T=366640 137600 0 0 $X=366350 $Y=137365
X1251 1 2 ICV_13 $T=366640 145440 1 0 $X=366350 $Y=141230
X1252 1 2 ICV_13 $T=366640 153280 0 0 $X=366350 $Y=153045
X1253 1 2 ICV_13 $T=366640 161120 0 0 $X=366350 $Y=160885
X1254 1 2 ICV_13 $T=371120 114080 0 0 $X=370830 $Y=113845
X1255 1 2 ICV_13 $T=371120 137600 1 0 $X=370830 $Y=133390
X1256 1 2 ICV_13 $T=382880 106240 0 0 $X=382590 $Y=106005
X1257 1 2 ICV_13 $T=408640 129760 1 0 $X=408350 $Y=125550
X1258 1 2 ICV_13 $T=408640 153280 0 0 $X=408350 $Y=153045
X1259 1 2 ICV_13 $T=417600 129760 1 0 $X=417310 $Y=125550
X1260 1 2 ICV_13 $T=418160 161120 1 0 $X=417870 $Y=156910
X1261 1 2 ICV_13 $T=429360 114080 0 0 $X=429070 $Y=113845
X1262 1 2 ICV_13 $T=429920 106240 0 0 $X=429630 $Y=106005
X1263 1 2 ICV_13 $T=450080 121920 0 0 $X=449790 $Y=121685
X1264 1 2 ICV_13 $T=450640 106240 0 0 $X=450350 $Y=106005
X1265 1 2 ICV_13 $T=459600 129760 1 0 $X=459310 $Y=125550
X1266 1 2 ICV_13 $T=470800 145440 1 0 $X=470510 $Y=141230
X1267 1 2 ICV_13 $T=470800 145440 0 0 $X=470510 $Y=145205
X1268 4 1 2 10 INVD1BWP7T $T=21680 168960 1 0 $X=21390 $Y=164750
X1269 8 1 2 913 INVD1BWP7T $T=23360 137600 1 0 $X=23070 $Y=133390
X1270 923 1 2 20 INVD1BWP7T $T=28400 153280 0 0 $X=28110 $Y=153045
X1271 917 1 2 43 INVD1BWP7T $T=38480 145440 1 0 $X=38190 $Y=141230
X1272 83 1 2 952 INVD1BWP7T $T=49680 145440 0 0 $X=49390 $Y=145205
X1273 75 1 2 954 INVD1BWP7T $T=50240 129760 1 0 $X=49950 $Y=125550
X1274 91 1 2 922 INVD1BWP7T $T=54720 114080 0 180 $X=52750 $Y=109870
X1275 932 1 2 97 INVD1BWP7T $T=54160 129760 1 0 $X=53870 $Y=125550
X1276 51 1 2 99 INVD1BWP7T $T=58640 114080 1 0 $X=58350 $Y=109870
X1277 48 1 2 116 INVD1BWP7T $T=58640 161120 0 0 $X=58350 $Y=160885
X1278 982 1 2 78 INVD1BWP7T $T=73200 129760 0 180 $X=71230 $Y=125550
X1279 163 1 2 971 INVD1BWP7T $T=87760 145440 0 180 $X=85790 $Y=141230
X1280 171 1 2 991 INVD1BWP7T $T=92240 129760 0 180 $X=90270 $Y=125550
X1281 207 1 2 1015 INVD1BWP7T $T=98960 114080 0 180 $X=96990 $Y=109870
X1282 211 1 2 1016 INVD1BWP7T $T=98960 121920 1 180 $X=96990 $Y=121685
X1283 242 1 2 221 INVD1BWP7T $T=110720 161120 0 180 $X=108750 $Y=156910
X1284 915 1 2 241 INVD1BWP7T $T=115200 161120 1 180 $X=113230 $Y=160885
X1285 272 1 2 1011 INVD1BWP7T $T=125840 153280 1 180 $X=123870 $Y=153045
X1286 1060 1 2 1062 INVD1BWP7T $T=131440 129760 0 0 $X=131150 $Y=129525
X1287 1072 1 2 1019 INVD1BWP7T $T=137600 161120 0 180 $X=135630 $Y=156910
X1288 1054 1 2 1094 INVD1BWP7T $T=143760 137600 0 180 $X=141790 $Y=133390
X1289 1061 1 2 315 INVD1BWP7T $T=143200 168960 1 0 $X=142910 $Y=164750
X1290 1101 1 2 1074 INVD1BWP7T $T=145440 137600 0 180 $X=143470 $Y=133390
X1291 1066 1 2 1099 INVD1BWP7T $T=151600 145440 0 180 $X=149630 $Y=141230
X1292 352 1 2 1119 INVD1BWP7T $T=166160 137600 0 180 $X=164190 $Y=133390
X1293 392 1 2 396 INVD1BWP7T $T=180160 168960 1 0 $X=179870 $Y=164750
X1294 390 1 2 378 INVD1BWP7T $T=183520 106240 0 0 $X=183230 $Y=106005
X1295 1163 1 2 458 INVD1BWP7T $T=222720 121920 1 0 $X=222430 $Y=117710
X1296 495 1 2 1209 INVD1BWP7T $T=259120 145440 0 0 $X=258830 $Y=145205
X1297 541 1 2 1251 INVD1BWP7T $T=293280 114080 0 180 $X=291310 $Y=109870
X1298 542 1 2 1258 INVD1BWP7T $T=292720 153280 0 0 $X=292430 $Y=153045
X1299 564 1 2 492 INVD1BWP7T $T=310080 168960 0 180 $X=308110 $Y=164750
X1300 594 1 2 1226 INVD1BWP7T $T=325200 161120 0 180 $X=323230 $Y=156910
X1301 680 1 2 678 INVD1BWP7T $T=392400 137600 0 180 $X=390430 $Y=133390
X1302 683 1 2 688 INVD1BWP7T $T=393520 161120 0 0 $X=393230 $Y=160885
X1303 1 2 ICV_14 $T=27840 114080 1 0 $X=27550 $Y=109870
X1304 1 2 ICV_14 $T=47440 114080 1 0 $X=47150 $Y=109870
X1305 1 2 ICV_14 $T=59760 161120 1 0 $X=59470 $Y=156910
X1306 1 2 ICV_14 $T=70400 161120 1 0 $X=70110 $Y=156910
X1307 1 2 ICV_14 $T=133120 168960 1 0 $X=132830 $Y=164750
X1308 1 2 ICV_14 $T=196400 121920 1 0 $X=196110 $Y=117710
X1309 1 2 ICV_14 $T=238400 153280 0 0 $X=238110 $Y=153045
X1310 1 2 ICV_14 $T=261920 106240 0 0 $X=261630 $Y=106005
X1311 1 2 ICV_14 $T=300560 129760 0 0 $X=300270 $Y=129525
X1312 1 2 ICV_14 $T=308960 161120 1 0 $X=308670 $Y=156910
X1313 1 2 ICV_14 $T=322400 153280 0 0 $X=322110 $Y=153045
X1314 1 2 ICV_14 $T=344240 137600 0 0 $X=343950 $Y=137365
X1315 1 2 ICV_14 $T=353760 137600 0 0 $X=353470 $Y=137365
X1316 1 2 ICV_14 $T=364400 114080 1 0 $X=364110 $Y=109870
X1317 1 2 ICV_14 $T=371120 129760 0 0 $X=370830 $Y=129525
X1318 1 2 ICV_14 $T=379520 129760 0 0 $X=379230 $Y=129525
X1319 1 2 ICV_14 $T=406400 114080 1 0 $X=406110 $Y=109870
X1320 486 503 1 2 BUFFD10BWP7T $T=251280 106240 0 0 $X=250990 $Y=106005
X1321 1009 201 1 2 BUFFD2BWP7T $T=95600 137600 0 0 $X=95310 $Y=137365
X1322 995 222 1 2 BUFFD2BWP7T $T=102320 137600 0 0 $X=102030 $Y=137365
X1323 990 244 1 2 BUFFD2BWP7T $T=107360 137600 0 0 $X=107070 $Y=137365
X1324 1012 313 1 2 BUFFD2BWP7T $T=142080 153280 0 0 $X=141790 $Y=153045
X1325 1013 314 1 2 BUFFD2BWP7T $T=142080 161120 1 0 $X=141790 $Y=156910
X1326 456 462 1 2 BUFFD2BWP7T $T=223280 145440 0 0 $X=222990 $Y=145205
X1327 1 2 DCAP16BWP7T $T=35120 161120 0 0 $X=34830 $Y=160885
X1328 1 2 DCAP16BWP7T $T=77120 129760 0 0 $X=76830 $Y=129525
X1329 1 2 DCAP16BWP7T $T=161120 121920 0 0 $X=160830 $Y=121685
X1330 1 2 DCAP16BWP7T $T=161120 129760 0 0 $X=160830 $Y=129525
X1331 1 2 DCAP16BWP7T $T=203120 129760 1 0 $X=202830 $Y=125550
X1332 1 2 DCAP16BWP7T $T=203120 161120 1 0 $X=202830 $Y=156910
X1333 1 2 DCAP16BWP7T $T=209840 168960 1 0 $X=209550 $Y=164750
X1334 1 2 DCAP16BWP7T $T=213200 137600 1 0 $X=212910 $Y=133390
X1335 1 2 DCAP16BWP7T $T=221040 129760 1 0 $X=220750 $Y=125550
X1336 1 2 DCAP16BWP7T $T=224400 121920 1 0 $X=224110 $Y=117710
X1337 1 2 DCAP16BWP7T $T=226080 168960 1 0 $X=225790 $Y=164750
X1338 1 2 DCAP16BWP7T $T=233360 114080 0 0 $X=233070 $Y=113845
X1339 1 2 DCAP16BWP7T $T=245120 153280 1 0 $X=244830 $Y=149070
X1340 1 2 DCAP16BWP7T $T=260800 145440 0 0 $X=260510 $Y=145205
X1341 1 2 DCAP16BWP7T $T=287120 161120 1 0 $X=286830 $Y=156910
X1342 1 2 DCAP16BWP7T $T=294960 121920 1 0 $X=294670 $Y=117710
X1343 1 2 DCAP16BWP7T $T=314000 145440 1 0 $X=313710 $Y=141230
X1344 1 2 DCAP16BWP7T $T=315120 121920 1 0 $X=314830 $Y=117710
X1345 1 2 DCAP16BWP7T $T=329120 145440 1 0 $X=328830 $Y=141230
X1346 1 2 DCAP16BWP7T $T=329120 153280 1 0 $X=328830 $Y=149070
X1347 1 2 DCAP16BWP7T $T=358240 121920 1 0 $X=357950 $Y=117710
X1348 1 2 DCAP16BWP7T $T=371120 121920 0 0 $X=370830 $Y=121685
X1349 1 2 DCAP16BWP7T $T=371120 137600 0 0 $X=370830 $Y=137365
X1350 1 2 DCAP16BWP7T $T=377280 114080 0 0 $X=376990 $Y=113845
X1351 1 2 DCAP16BWP7T $T=383440 114080 1 0 $X=383150 $Y=109870
X1352 1 2 DCAP16BWP7T $T=389040 153280 0 0 $X=388750 $Y=153045
X1353 1 2 DCAP16BWP7T $T=402480 145440 1 0 $X=402190 $Y=141230
X1354 1 2 DCAP16BWP7T $T=422640 129760 1 0 $X=422350 $Y=125550
X1355 1 2 DCAP16BWP7T $T=424320 145440 0 0 $X=424030 $Y=145205
X1356 1 2 DCAP16BWP7T $T=430480 161120 0 0 $X=430190 $Y=160885
X1357 1 2 DCAP16BWP7T $T=443360 121920 1 0 $X=443070 $Y=117710
X1358 1 2 DCAP16BWP7T $T=443360 145440 1 0 $X=443070 $Y=141230
X1359 1 2 DCAP16BWP7T $T=445040 153280 0 0 $X=444750 $Y=153045
X1360 1 2 DCAP16BWP7T $T=455120 137600 1 0 $X=454830 $Y=133390
X1361 949 1 2 76 CKND1BWP7T $T=50240 168960 0 180 $X=48270 $Y=164750
X1362 95 1 2 88 CKND1BWP7T $T=54160 161120 0 180 $X=52190 $Y=156910
X1363 238 1 2 1036 CKND1BWP7T $T=130320 153280 0 180 $X=128350 $Y=149070
X1364 537 1 2 1243 CKND1BWP7T $T=289920 161120 0 0 $X=289630 $Y=160885
X1365 604 1 2 610 CKND1BWP7T $T=348160 161120 0 180 $X=346190 $Y=156910
X1366 1144 1 2 1312 CKND1BWP7T $T=359360 114080 0 180 $X=357390 $Y=109870
X1367 676 1 2 1333 CKND1BWP7T $T=387920 153280 0 180 $X=385950 $Y=149070
X1368 619 1 2 1373 CKND1BWP7T $T=406400 145440 0 0 $X=406110 $Y=145205
X1369 717 1 2 712 CKND1BWP7T $T=420400 114080 0 180 $X=418430 $Y=109870
X1370 718 1 2 700 CKND1BWP7T $T=420400 114080 1 0 $X=420110 $Y=109870
X1371 102 130 1 2 INVD4BWP7T $T=65360 153280 0 0 $X=65070 $Y=153045
X1372 486 1 2 480 BUFFD3BWP7T $T=237280 121920 0 180 $X=233070 $Y=117710
X1373 674 1345 238 1 2 CKXOR2D4BWP7T $T=388480 161120 0 180 $X=375870 $Y=156910
X1374 1238 421 2 1241 1 527 1220 AOI22D1BWP7T $T=279840 121920 0 180 $X=275630 $Y=117710
X1375 1214 421 2 1229 1 527 1246 AOI22D1BWP7T $T=277600 129760 1 0 $X=277310 $Y=125550
X1376 613 611 2 608 1 1293 601 AOI22D1BWP7T $T=340320 168960 0 180 $X=336110 $Y=164750
X1377 1309 1187 2 626 1 628 1314 AOI22D1BWP7T $T=347600 137600 1 0 $X=347310 $Y=133390
X1378 622 1312 2 629 1 1144 1317 AOI22D1BWP7T $T=348720 114080 1 0 $X=348430 $Y=109870
X1379 1313 1187 2 1311 1 628 1305 AOI22D1BWP7T $T=349840 137600 0 0 $X=349550 $Y=137365
X1380 643 1312 2 1326 1 1144 1330 AOI22D1BWP7T $T=363280 114080 1 180 $X=359070 $Y=113845
X1381 1355 666 2 1344 1 662 1325 AOI22D1BWP7T $T=382320 161120 1 180 $X=378110 $Y=160885
X1382 661 1312 2 664 1 1321 1341 AOI22D1BWP7T $T=378960 106240 0 0 $X=378670 $Y=106005
X1383 1352 1312 2 665 1 1321 1343 AOI22D1BWP7T $T=383440 114080 0 180 $X=379230 $Y=109870
X1384 1351 666 2 667 1 662 1338 AOI22D1BWP7T $T=384560 137600 1 180 $X=380350 $Y=137365
X1385 1356 685 2 684 1 462 1361 AOI22D1BWP7T $T=392960 129760 0 0 $X=392670 $Y=129525
X1386 695 685 2 697 1 462 1364 AOI22D1BWP7T $T=399680 145440 0 0 $X=399390 $Y=145205
X1387 580 2 374 1 CKND12BWP7T $T=313440 121920 0 0 $X=313150 $Y=121685
X1388 1181 476 1 2 BUFFD8BWP7T $T=227200 129760 0 0 $X=226910 $Y=129525
X1389 1173 477 1 2 BUFFD8BWP7T $T=240080 129760 0 180 $X=230830 $Y=125550
X1390 578 561 1 2 BUFFD8BWP7T $T=315120 121920 0 180 $X=305870 $Y=117710
X1391 605 525 1 2 BUFFD8BWP7T $T=336960 129760 0 0 $X=336670 $Y=129525
X1392 437 578 1 2 BUFFD8BWP7T $T=417600 129760 0 0 $X=417310 $Y=129525
X1393 1178 455 1 2 BUFFD6BWP7T $T=219360 168960 1 0 $X=219070 $Y=164750
X1394 28 22 2 1 INVD2BWP7T $T=27840 114080 0 180 $X=25310 $Y=109870
X1395 939 45 2 1 INVD2BWP7T $T=44640 129760 0 180 $X=42110 $Y=125550
X1396 127 79 2 1 INVD2BWP7T $T=63120 161120 1 180 $X=60590 $Y=160885
X1397 973 149 2 1 INVD2BWP7T $T=69840 137600 0 0 $X=69550 $Y=137365
X1398 169 984 2 1 INVD2BWP7T $T=86080 145440 0 180 $X=83550 $Y=141230
X1399 175 930 2 1 INVD2BWP7T $T=95040 145440 0 180 $X=92510 $Y=141230
X1400 182 256 2 1 INVD2BWP7T $T=130880 161120 1 180 $X=128350 $Y=160885
X1401 1147 408 2 1 INVD2BWP7T $T=189120 129760 1 180 $X=186590 $Y=129525
X1402 459 1191 2 1 INVD2BWP7T $T=224400 153280 1 0 $X=224110 $Y=149070
X1403 494 1242 2 1 INVD2BWP7T $T=279840 137600 0 0 $X=279550 $Y=137365
X1404 538 1254 2 1 INVD2BWP7T $T=290480 153280 0 0 $X=290190 $Y=153045
X1405 624 655 2 1 INVD2BWP7T $T=376720 137600 0 180 $X=374190 $Y=133390
X1406 1381 771 2 1 INVD2BWP7T $T=458480 161120 0 0 $X=458190 $Y=160885
X1407 1280 774 2 1 INVD2BWP7T $T=460720 114080 1 0 $X=460430 $Y=109870
X1408 1384 781 2 1 INVD2BWP7T $T=462960 114080 1 0 $X=462670 $Y=109870
X1409 1385 782 2 1 INVD2BWP7T $T=463520 129760 1 0 $X=463230 $Y=125550
X1410 788 785 2 1 INVD2BWP7T $T=466880 137600 0 180 $X=464350 $Y=133390
X1411 793 796 2 1 INVD2BWP7T $T=469120 121920 1 0 $X=468830 $Y=117710
X1412 794 797 2 1 INVD2BWP7T $T=469680 114080 1 0 $X=469390 $Y=109870
X1413 1387 800 2 1 INVD2BWP7T $T=471920 114080 1 0 $X=471630 $Y=109870
X1414 1190 1168 1 2 1193 CKXOR2D1BWP7T $T=223840 161120 0 0 $X=223550 $Y=160885
X1415 1225 1209 1 2 1219 CKXOR2D1BWP7T $T=266960 145440 0 180 $X=261630 $Y=141230
X1416 495 1265 1 2 1264 CKXOR2D1BWP7T $T=296080 145440 0 0 $X=295790 $Y=145205
X1417 1248 553 1 2 539 CKXOR2D1BWP7T $T=297200 168960 1 0 $X=296910 $Y=164750
X1418 1264 551 1 2 1263 CKXOR2D1BWP7T $T=302800 161120 0 180 $X=297470 $Y=156910
X1419 1144 522 1 2 582 CKXOR2D1BWP7T $T=310640 114080 0 0 $X=310350 $Y=113845
X1420 583 1144 1 2 1288 CKXOR2D1BWP7T $T=317360 114080 1 0 $X=317070 $Y=109870
X1421 1277 591 1 2 1283 CKXOR2D1BWP7T $T=319600 137600 0 0 $X=319310 $Y=137365
X1422 1288 584 1 2 1285 CKXOR2D1BWP7T $T=320160 137600 1 0 $X=319870 $Y=133390
X1423 603 616 1 2 1300 CKXOR2D1BWP7T $T=339200 137600 0 0 $X=338910 $Y=137365
X1424 462 635 1 2 1366 CKXOR2D1BWP7T $T=396320 121920 1 0 $X=396030 $Y=117710
X1425 494 1200 1072 1 2 CKXOR2D2BWP7T $T=241200 137600 0 180 $X=234750 $Y=133390
X1426 505 497 1105 1 2 CKXOR2D2BWP7T $T=254080 145440 0 180 $X=247630 $Y=141230
X1427 1298 619 927 1 2 CKXOR2D2BWP7T $T=348160 153280 0 180 $X=341710 $Y=149070
X1428 624 1304 618 1 2 CKXOR2D2BWP7T $T=349840 121920 0 180 $X=343390 $Y=117710
X1429 722 1370 1023 1 2 CKXOR2D2BWP7T $T=424320 145440 1 180 $X=417870 $Y=145205
X1430 2 1 DCAP32BWP7T $T=329120 121920 0 0 $X=328830 $Y=121685
X1431 2 1 DCAP32BWP7T $T=371120 153280 0 0 $X=370830 $Y=153045
X1432 2 1 DCAP32BWP7T $T=392400 137600 1 0 $X=392110 $Y=133390
X1433 2 1 DCAP32BWP7T $T=455120 106240 0 0 $X=454830 $Y=106005
X1434 2 1 DCAP32BWP7T $T=455120 114080 0 0 $X=454830 $Y=113845
X1435 2 1 DCAP32BWP7T $T=455120 161120 1 0 $X=454830 $Y=156910
X1436 263 1067 1033 1062 1 2 OAI21D0BWP7T $T=125280 114080 0 0 $X=124990 $Y=113845
X1437 1223 1230 517 477 1 2 OAI21D0BWP7T $T=270320 121920 1 0 $X=270030 $Y=117710
X1438 1249 1261 544 477 1 2 OAI21D0BWP7T $T=294960 129760 1 0 $X=294670 $Y=125550
X1439 620 1303 621 1173 1 2 OAI21D0BWP7T $T=347040 114080 1 180 $X=343950 $Y=113845
X1440 1319 1329 641 477 1 2 OAI21D0BWP7T $T=360480 145440 1 0 $X=360190 $Y=141230
X1441 652 653 656 477 1 2 OAI21D0BWP7T $T=373920 106240 0 0 $X=373630 $Y=106005
X1442 1330 1332 657 1337 1 2 OAI21D0BWP7T $T=374480 114080 0 0 $X=374190 $Y=113845
X1443 1334 1339 658 485 1 2 OAI21D0BWP7T $T=376720 129760 0 0 $X=376430 $Y=129525
X1444 1314 1335 649 485 1 2 OAI21D0BWP7T $T=377840 145440 0 0 $X=377550 $Y=145205
X1445 1338 1346 663 485 1 2 OAI21D0BWP7T $T=381760 153280 1 0 $X=381470 $Y=149070
X1446 1343 1349 673 1353 1 2 OAI21D0BWP7T $T=384560 121920 1 0 $X=384270 $Y=117710
X1447 1348 1350 670 485 1 2 OAI21D0BWP7T $T=385120 129760 0 0 $X=384830 $Y=129525
X1448 1375 1374 696 1365 1 2 OAI21D0BWP7T $T=405280 129760 1 180 $X=402190 $Y=129525
X1449 1379 1378 710 485 1 2 OAI21D0BWP7T $T=422080 114080 0 0 $X=421790 $Y=113845
X1450 546 1219 547 1 2 1266 MUX2ND1BWP7T $T=293840 161120 0 0 $X=293550 $Y=160885
X1451 452 1168 1 2 1189 XNR2D1BWP7T $T=219920 153280 0 0 $X=219630 $Y=153045
X1452 1193 492 1 2 1203 XNR2D1BWP7T $T=235600 161120 0 0 $X=235310 $Y=160885
X1453 1224 1184 1 2 528 XNR2D1BWP7T $T=272000 153280 0 0 $X=271710 $Y=153045
X1454 1237 1184 1 2 1248 XNR2D1BWP7T $T=276480 168960 1 0 $X=276190 $Y=164750
X1455 581 1165 1 2 1277 XNR2D1BWP7T $T=316800 137600 0 180 $X=311470 $Y=133390
X1456 589 1279 1 2 1273 XNR2D1BWP7T $T=322400 153280 1 180 $X=317070 $Y=153045
X1457 25 24 2 1 CKND2BWP7T $T=26720 161120 0 180 $X=24190 $Y=156910
X1458 12 916 2 1 CKND2BWP7T $T=31200 137600 1 180 $X=28670 $Y=137365
X1459 475 511 2 1 CKND2BWP7T $T=256320 145440 1 0 $X=256030 $Y=141230
X1460 1302 769 2 1 CKND2BWP7T $T=457920 121920 1 0 $X=457630 $Y=117710
X1461 929 1 2 52 CKND0BWP7T $T=39040 114080 1 0 $X=38750 $Y=109870
X1462 195 1 2 1001 CKND0BWP7T $T=96160 137600 0 180 $X=94190 $Y=133390
X1463 229 1 2 217 CKND0BWP7T $T=107360 161120 0 180 $X=105390 $Y=156910
X1464 1042 1 2 1051 CKND0BWP7T $T=122480 145440 0 0 $X=122190 $Y=145205
X1465 332 1 2 1117 CKND0BWP7T $T=153280 145440 1 180 $X=151310 $Y=145205
X1466 595 1 2 598 CKND0BWP7T $T=331920 106240 0 0 $X=331630 $Y=106005
X1467 714 1 2 711 CKND0BWP7T $T=419840 137600 0 180 $X=417870 $Y=133390
X1468 371 2 401 1135 388 326 1 AOI22D2BWP7T $T=184640 145440 0 180 $X=177630 $Y=141230
X1469 501 2 1209 1198 495 1207 1 AOI22D2BWP7T $T=255760 145440 1 180 $X=248750 $Y=145205
X1470 507 2 1209 496 495 498 1 AOI22D2BWP7T $T=255760 168960 0 180 $X=248750 $Y=164750
X1471 1269 2 1183 568 563 548 1 AOI22D2BWP7T $T=302800 129760 1 0 $X=302510 $Y=125550
X1472 573 2 1183 562 563 1276 1 AOI22D2BWP7T $T=312880 129760 1 180 $X=305870 $Y=129525
X1473 1189 473 1194 1197 1 2 MUX2ND0BWP7T $T=229440 161120 1 0 $X=229150 $Y=156910
X1474 1273 585 587 1287 1 2 MUX2ND0BWP7T $T=316800 161120 0 0 $X=316510 $Y=160885
X1475 593 604 610 1296 1 2 MUX2ND0BWP7T $T=335280 121920 1 0 $X=334990 $Y=117710
X1476 945 968 966 78 960 2 1 AOI22D0BWP7T $T=62560 129760 1 180 $X=58910 $Y=129525
X1477 1168 1192 466 470 1189 2 1 AOI22D0BWP7T $T=227200 153280 0 0 $X=226910 $Y=153045
X1478 1203 1202 1193 485 482 2 1 AOI22D0BWP7T $T=238960 161120 0 180 $X=235310 $Y=156910
X1479 1043 1 2 1058 CKBD0BWP7T $T=121920 129760 1 0 $X=121630 $Y=125550
X1480 266 1 2 1109 CKBD0BWP7T $T=147120 114080 1 0 $X=146830 $Y=109870
X1481 1151 1 2 1171 CKBD0BWP7T $T=214880 153280 1 0 $X=214590 $Y=149070
X1482 1165 1 2 1279 CKBD0BWP7T $T=310640 153280 0 0 $X=310350 $Y=153045
X1483 1364 1 2 1375 CKBD0BWP7T $T=405840 129760 0 0 $X=405550 $Y=129525
X1484 378 391 393 394 2 1 397 AO211D1BWP7T $T=179040 106240 0 0 $X=178750 $Y=106005
X1485 913 2 914 3 1 NR2D1BWP7T $T=28960 137600 0 180 $X=26430 $Y=133390
X1486 933 2 46 927 1 NR2D1BWP7T $T=41840 137600 0 180 $X=39310 $Y=133390
X1487 939 2 932 62 1 NR2D1BWP7T $T=44640 129760 1 0 $X=44350 $Y=125550
X1488 99 2 957 90 1 NR2D1BWP7T $T=56400 106240 1 180 $X=53870 $Y=106005
X1489 101 2 969 125 1 NR2D1BWP7T $T=73200 121920 1 180 $X=70670 $Y=121685
X1490 930 2 198 915 1 NR2D1BWP7T $T=95040 161120 0 0 $X=94750 $Y=160885
X1491 1022 2 203 1011 1 NR2D1BWP7T $T=99520 161120 1 180 $X=96990 $Y=160885
X1492 234 2 246 1039 1 NR2D1BWP7T $T=109600 114080 0 0 $X=109310 $Y=113845
X1493 163 2 1041 1023 1 NR2D1BWP7T $T=124160 153280 1 180 $X=121630 $Y=153045
X1494 1070 2 279 1039 1 NR2D1BWP7T $T=130880 121920 0 180 $X=128350 $Y=117710
X1495 182 2 286 1072 1 NR2D1BWP7T $T=130880 168960 1 0 $X=130590 $Y=164750
X1496 1036 2 1077 1072 1 NR2D1BWP7T $T=133120 161120 0 0 $X=132830 $Y=160885
X1497 293 2 1063 1031 1 NR2D1BWP7T $T=135920 137600 0 180 $X=133390 $Y=133390
X1498 208 2 1071 301 1 NR2D1BWP7T $T=135920 106240 0 0 $X=135630 $Y=106005
X1499 366 2 354 362 1 NR2D1BWP7T $T=170080 168960 0 180 $X=167550 $Y=164750
X1500 326 2 1136 381 1 NR2D1BWP7T $T=182400 129760 1 180 $X=179870 $Y=129525
X1501 357 2 1149 381 1 NR2D1BWP7T $T=196400 153280 1 0 $X=196110 $Y=149070
X1502 430 2 427 1162 1 NR2D1BWP7T $T=205920 114080 0 0 $X=205630 $Y=113845
X1503 1198 2 1201 478 1 NR2D1BWP7T $T=238960 145440 1 180 $X=236430 $Y=145205
X1504 495 2 1199 499 1 NR2D1BWP7T $T=248480 161120 1 0 $X=248190 $Y=156910
X1505 48 934 930 25 1 2 AOI21D0BWP7T $T=41280 153280 1 180 $X=38190 $Y=153045
X1506 156 993 78 997 1 2 AOI21D0BWP7T $T=80480 121920 1 0 $X=80190 $Y=117710
X1507 988 1002 173 174 1 2 AOI21D0BWP7T $T=85520 106240 0 0 $X=85230 $Y=106005
X1508 330 1113 1027 1066 1 2 AOI21D0BWP7T $T=148800 129760 1 0 $X=148510 $Y=125550
X1509 1118 1115 338 1094 1 2 AOI21D0BWP7T $T=153280 114080 1 180 $X=150190 $Y=113845
X1510 1158 1150 427 1146 1 2 AOI21D0BWP7T $T=199200 114080 1 180 $X=196110 $Y=113845
X1511 438 1160 434 390 1 2 AOI21D0BWP7T $T=209280 106240 1 180 $X=206190 $Y=106005
X1512 1223 1228 517 1230 1 2 AOI21D0BWP7T $T=265840 114080 0 0 $X=265550 $Y=113845
X1513 532 1247 530 529 1 2 AOI21D0BWP7T $T=282640 106240 1 180 $X=279550 $Y=106005
X1514 1249 1253 544 1261 1 2 AOI21D0BWP7T $T=292160 121920 1 0 $X=291870 $Y=117710
X1515 1287 1271 477 1281 1 2 AOI21D0BWP7T $T=318480 145440 1 180 $X=315390 $Y=145205
X1516 1319 1322 641 1329 1 2 AOI21D0BWP7T $T=359360 137600 0 0 $X=359070 $Y=137365
X1517 1314 1324 649 1335 1 2 AOI21D0BWP7T $T=363840 145440 1 0 $X=363550 $Y=141230
X1518 1334 1336 658 1339 1 2 AOI21D0BWP7T $T=374480 129760 1 0 $X=374190 $Y=125550
X1519 1330 1337 657 484 1 2 AOI21D0BWP7T $T=375600 121920 1 0 $X=375310 $Y=117710
X1520 1338 1340 663 1346 1 2 AOI21D0BWP7T $T=378960 153280 1 0 $X=378670 $Y=149070
X1521 1348 1347 670 1350 1 2 AOI21D0BWP7T $T=381760 137600 1 0 $X=381470 $Y=133390
X1522 654 659 672 675 1 2 AOI21D0BWP7T $T=384560 168960 1 0 $X=384270 $Y=164750
X1523 1343 1353 673 484 1 2 AOI21D0BWP7T $T=387360 121920 1 0 $X=387070 $Y=117710
X1524 1364 1365 696 484 1 2 AOI21D0BWP7T $T=399120 129760 0 0 $X=398830 $Y=129525
X1525 1379 1376 710 1378 1 2 AOI21D0BWP7T $T=419840 114080 1 180 $X=416750 $Y=113845
X1526 926 34 922 30 2 1 33 NR4D1BWP7T $T=31200 106240 1 180 $X=25310 $Y=106005
X1527 974 947 131 125 2 1 123 NR4D1BWP7T $T=67040 121920 1 180 $X=61150 $Y=121685
X1528 977 140 947 137 2 1 963 NR4D1BWP7T $T=69840 121920 0 180 $X=63950 $Y=117710
X1529 1024 1016 189 1014 2 1 206 NR4D1BWP7T $T=101760 121920 0 180 $X=95870 $Y=117710
X1530 1032 234 228 1021 2 1 190 NR4D1BWP7T $T=109040 114080 1 180 $X=103150 $Y=113845
X1531 276 258 269 1047 2 1 260 NR4D1BWP7T $T=127520 114080 0 180 $X=121630 $Y=109870
X1532 1064 281 1015 287 2 1 288 NR4D1BWP7T $T=128640 114080 1 0 $X=128350 $Y=109870
X1533 1069 1075 290 284 2 1 282 NR4D1BWP7T $T=135360 121920 1 180 $X=129470 $Y=121685
X1534 1079 1070 239 298 2 1 297 NR4D1BWP7T $T=132000 114080 0 0 $X=131710 $Y=113845
X1535 1095 1086 306 1034 2 1 291 NR4D1BWP7T $T=140960 121920 0 180 $X=135070 $Y=117710
X1536 1091 318 311 310 2 1 309 NR4D1BWP7T $T=147120 114080 0 180 $X=141230 $Y=109870
X1537 1122 208 358 363 2 1 361 NR4D1BWP7T $T=164480 106240 0 0 $X=164190 $Y=106005
X1538 1154 1138 1149 413 2 1 416 NR4D1BWP7T $T=195280 153280 1 180 $X=189390 $Y=153045
X1539 434 463 465 471 2 1 467 NR4D1BWP7T $T=226080 106240 0 0 $X=225790 $Y=106005
X1540 1177 460 463 490 2 1 487 NR4D1BWP7T $T=233920 106240 0 0 $X=233630 $Y=106005
X1541 39 2 58 44 53 13 1 AOI31D2BWP7T $T=37920 121920 1 0 $X=37630 $Y=117710
X1542 1066 2 1083 1068 1045 1079 1 AOI31D2BWP7T $T=129760 145440 1 0 $X=129470 $Y=141230
X1543 1138 2 1145 368 350 326 1 AOI31D2BWP7T $T=184080 145440 0 0 $X=183790 $Y=145205
X1544 423 420 419 1148 2 1 1147 OR4D1BWP7T $T=195280 114080 0 180 $X=190510 $Y=109870
X1545 927 44 19 59 1 2 944 OA31D0BWP7T $T=42960 137600 1 0 $X=42670 $Y=133390
X1546 964 135 138 78 1 2 980 OA31D0BWP7T $T=65360 129760 1 0 $X=65070 $Y=125550
X1547 68 126 162 966 1 2 999 OA31D0BWP7T $T=80480 114080 0 0 $X=80190 $Y=113845
X1548 981 2 141 24 130 1 AOI21D2BWP7T $T=70400 161120 0 180 $X=65070 $Y=156910
X1549 1011 2 196 57 984 1 AOI21D2BWP7T $T=96160 153280 0 180 $X=90830 $Y=149070
X1550 1060 2 1076 1063 1048 1 AOI21D2BWP7T $T=138720 145440 1 180 $X=133390 $Y=145205
X1551 1094 2 1087 1082 1091 1 AOI21D2BWP7T $T=143760 145440 0 180 $X=138430 $Y=141230
X1552 1074 2 1106 1085 1110 1 AOI21D2BWP7T $T=144320 145440 1 0 $X=144030 $Y=141230
X1553 1119 2 331 328 326 1 AOI21D2BWP7T $T=152160 161120 1 180 $X=146830 $Y=160885
X1554 372 2 379 378 377 1 AOI21D2BWP7T $T=170640 106240 0 0 $X=170350 $Y=106005
X1555 390 2 1134 384 383 1 AOI21D2BWP7T $T=180160 114080 0 180 $X=174830 $Y=109870
X1556 388 2 1133 386 389 1 AOI21D2BWP7T $T=180720 145440 1 180 $X=175390 $Y=145205
X1557 337 2 1143 328 336 1 AOI21D2BWP7T $T=190800 153280 1 0 $X=190510 $Y=149070
X1558 3 1 9 12 2 ND2D1BWP7T $T=21680 137600 0 0 $X=21390 $Y=137365
X1559 15 1 17 12 2 ND2D1BWP7T $T=25600 114080 0 180 $X=23070 $Y=109870
X1560 20 1 26 24 2 ND2D1BWP7T $T=24480 168960 1 0 $X=24190 $Y=164750
X1561 916 1 27 914 2 ND2D1BWP7T $T=27280 121920 0 180 $X=24750 $Y=117710
X1562 913 1 16 3 2 ND2D1BWP7T $T=28960 137600 1 0 $X=28670 $Y=133390
X1563 15 1 42 45 2 ND2D1BWP7T $T=38480 106240 0 0 $X=38190 $Y=106005
X1564 44 1 917 928 2 ND2D1BWP7T $T=42400 145440 0 180 $X=39870 $Y=141230
X1565 36 1 51 23 2 ND2D1BWP7T $T=40720 106240 0 0 $X=40430 $Y=106005
X1566 5 1 937 55 2 ND2D1BWP7T $T=41840 114080 0 0 $X=41550 $Y=113845
X1567 43 1 939 13 2 ND2D1BWP7T $T=45760 145440 0 180 $X=43230 $Y=141230
X1568 69 1 924 56 2 ND2D1BWP7T $T=46320 114080 1 180 $X=43790 $Y=113845
X1569 63 1 941 51 2 ND2D1BWP7T $T=45760 106240 0 0 $X=45470 $Y=106005
X1570 72 1 935 80 2 ND2D1BWP7T $T=48000 106240 0 0 $X=47710 $Y=106005
X1571 954 1 947 94 2 ND2D1BWP7T $T=51920 121920 1 0 $X=51630 $Y=117710
X1572 109 1 946 106 2 ND2D1BWP7T $T=59760 161120 0 180 $X=57230 $Y=156910
X1573 130 1 106 124 2 ND2D1BWP7T $T=64240 168960 0 180 $X=61710 $Y=164750
X1574 116 1 146 143 2 ND2D1BWP7T $T=67600 168960 1 0 $X=67310 $Y=164750
X1575 130 1 127 153 2 ND2D1BWP7T $T=69280 153280 0 0 $X=68990 $Y=153045
X1576 1001 1 982 176 2 ND2D1BWP7T $T=90560 129760 1 180 $X=88030 $Y=129525
X1577 194 1 190 187 2 ND2D1BWP7T $T=94480 114080 0 180 $X=91950 $Y=109870
X1578 176 1 133 195 2 ND2D1BWP7T $T=92240 137600 1 0 $X=91950 $Y=133390
X1579 213 1 1025 212 2 ND2D1BWP7T $T=101200 106240 0 0 $X=100910 $Y=106005
X1580 971 1 1022 1023 2 ND2D1BWP7T $T=101760 145440 0 0 $X=101470 $Y=145205
X1581 1023 1 159 221 2 ND2D1BWP7T $T=105120 153280 0 0 $X=104830 $Y=153045
X1582 245 1 1031 1020 2 ND2D1BWP7T $T=109600 137600 0 180 $X=107070 $Y=133390
X1583 1036 1 973 229 2 ND2D1BWP7T $T=110160 145440 1 180 $X=107630 $Y=145205
X1584 256 1 252 1042 2 ND2D1BWP7T $T=115200 168960 0 180 $X=112670 $Y=164750
X1585 240 1 1047 251 2 ND2D1BWP7T $T=121920 121920 1 0 $X=121630 $Y=117710
X1586 265 1 1055 1049 2 ND2D1BWP7T $T=123600 106240 0 0 $X=123310 $Y=106005
X1587 1072 1 938 238 2 ND2D1BWP7T $T=133120 161120 1 180 $X=130590 $Y=160885
X1588 1071 1 1075 1052 2 ND2D1BWP7T $T=132560 129760 1 0 $X=132270 $Y=125550
X1589 299 1 300 1077 2 ND2D1BWP7T $T=138720 161120 1 180 $X=136190 $Y=160885
X1590 251 1 1086 316 2 ND2D1BWP7T $T=143200 121920 1 0 $X=142910 $Y=117710
X1591 213 1 320 280 2 ND2D1BWP7T $T=144880 106240 0 0 $X=144590 $Y=106005
X1592 332 1 1060 1105 2 ND2D1BWP7T $T=149360 145440 1 180 $X=146830 $Y=145205
X1593 1105 1 1066 1117 2 ND2D1BWP7T $T=149360 145440 0 0 $X=149070 $Y=145205
X1594 375 1 371 353 2 ND2D1BWP7T $T=172320 168960 0 180 $X=169790 $Y=164750
X1595 356 1 1128 1131 2 ND2D1BWP7T $T=170640 161120 1 0 $X=170350 $Y=156910
X1596 417 1 352 399 2 ND2D1BWP7T $T=190240 161120 0 180 $X=187710 $Y=156910
X1597 430 1 390 1162 2 ND2D1BWP7T $T=210400 114080 1 180 $X=207870 $Y=113845
X1598 421 1 1222 446 2 ND2D1BWP7T $T=279280 145440 0 0 $X=278990 $Y=145205
X1599 1279 1 559 446 2 ND2D1BWP7T $T=316800 161120 0 180 $X=314270 $Y=156910
X1600 127 1 106 952 2 950 930 OAI211D1BWP7T $T=64240 153280 1 180 $X=60590 $Y=153045
X1601 967 1 968 128 2 948 133 OAI211D1BWP7T $T=61440 137600 1 0 $X=61150 $Y=133390
X1602 976 1 151 926 2 990 991 OAI211D1BWP7T $T=69840 129760 0 0 $X=69550 $Y=129525
X1603 970 1 993 168 2 1003 133 OAI211D1BWP7T $T=83280 121920 1 0 $X=82990 $Y=117710
X1604 178 1 1002 184 2 1008 991 OAI211D1BWP7T $T=88320 106240 0 0 $X=88030 $Y=106005
X1605 1018 1 157 4 2 224 1022 OAI211D1BWP7T $T=105680 161120 1 180 $X=102030 $Y=160885
X1606 1050 1 1067 1069 2 1073 1074 OAI211D1BWP7T $T=130320 137600 1 0 $X=130030 $Y=133390
X1607 1104 1 1084 312 2 1093 1060 OAI211D1BWP7T $T=146560 129760 1 180 $X=142910 $Y=129525
X1608 403 1 409 410 2 1146 412 OAI211D1BWP7T $T=186880 106240 0 0 $X=186590 $Y=106005
X1609 1151 1 1145 388 2 1174 385 OAI211D1BWP7T $T=213760 153280 0 0 $X=213470 $Y=153045
X1610 1202 1 1192 484 2 489 1197 OAI211D1BWP7T $T=238400 153280 1 180 $X=234750 $Y=153045
X1611 1222 1 1221 1220 2 1200 1195 OAI211D1BWP7T $T=264720 121920 0 180 $X=261070 $Y=117710
X1612 1222 1 1245 1246 2 535 1195 OAI211D1BWP7T $T=279840 121920 1 0 $X=279550 $Y=117710
X1613 559 1 1271 1273 2 566 1195 OAI211D1BWP7T $T=305600 145440 0 0 $X=305310 $Y=145205
X1614 531 1 1308 1305 2 1304 1195 OAI211D1BWP7T $T=347600 145440 0 180 $X=343950 $Y=141230
X1615 1332 1 1331 1317 2 642 545 OAI211D1BWP7T $T=364400 114080 0 180 $X=360750 $Y=109870
X1616 1349 1 1342 1341 2 1345 545 OAI211D1BWP7T $T=381200 129760 0 180 $X=377550 $Y=125550
X1617 1374 1 1372 1361 2 1370 545 OAI211D1BWP7T $T=404720 121920 1 180 $X=401070 $Y=121685
X1618 67 2 936 32 98 1 104 NR4D2BWP7T $T=44640 161120 0 0 $X=44350 $Y=160885
X1619 1017 2 210 1026 208 1 1027 NR4D2BWP7T $T=95040 129760 0 0 $X=94750 $Y=129525
X1620 481 2 465 469 460 1 472 NR4D2BWP7T $T=236720 114080 0 180 $X=223550 $Y=109870
X1621 915 2 48 158 1 NR2XD0BWP7T $T=82160 168960 0 180 $X=79630 $Y=164750
X1622 218 1 216 207 212 1017 2 ND4D1BWP7T $T=103440 114080 0 180 $X=99230 $Y=109870
X1623 231 1 240 236 226 1038 2 ND4D1BWP7T $T=106800 121920 0 0 $X=106510 $Y=121685
X1624 275 1 277 1049 280 1065 2 ND4D1BWP7T $T=126960 106240 0 0 $X=126670 $Y=106005
X1625 89 951 955 84 78 1 2 OAI31D1BWP7T $T=53600 137600 0 180 $X=49390 $Y=133390
X1626 959 117 967 111 105 1 2 OAI31D1BWP7T $T=61440 121920 1 180 $X=57230 $Y=121685
X1627 129 114 970 122 105 1 2 OAI31D1BWP7T $T=64240 114080 1 180 $X=60030 $Y=113845
X1628 113 131 996 161 966 1 2 OAI31D1BWP7T $T=79920 114080 1 0 $X=79630 $Y=109870
X1629 163 221 1005 217 215 1 2 OAI31D1BWP7T $T=105120 153280 1 180 $X=100910 $Y=153045
X1630 1038 259 1050 268 1054 1 2 OAI31D1BWP7T $T=121920 137600 1 0 $X=121630 $Y=133390
X1631 1046 1055 1059 1028 1062 1 2 OAI31D1BWP7T $T=124720 121920 0 0 $X=124430 $Y=121685
X1632 1038 255 1084 303 1054 1 2 OAI31D1BWP7T $T=136480 129760 0 0 $X=136190 $Y=129525
X1633 302 261 1088 1090 1054 1 2 OAI31D1BWP7T $T=138160 121920 0 0 $X=137870 $Y=121685
X1634 255 311 1103 323 1101 1 2 OAI31D1BWP7T $T=145440 121920 1 0 $X=145150 $Y=117710
X1635 260 290 1112 347 1099 1 2 OAI31D1BWP7T $T=153280 121920 0 0 $X=152990 $Y=121685
X1636 975 958 147 987 982 1 2 AOI31D0BWP7T $T=68720 114080 0 0 $X=68430 $Y=113845
X1637 983 150 96 989 154 1 2 AOI31D0BWP7T $T=69840 121920 1 0 $X=69550 $Y=117710
X1638 1044 1063 279 1057 1074 1 2 AOI31D0BWP7T $T=126960 137600 0 0 $X=126670 $Y=137365
X1639 1078 304 305 1089 1074 1 2 AOI31D0BWP7T $T=138160 114080 1 0 $X=137870 $Y=109870
X1640 321 1081 1068 1102 1074 1 2 AOI31D0BWP7T $T=146560 129760 0 180 $X=142910 $Y=125550
X1641 1032 1109 335 1116 1066 1 2 AOI31D0BWP7T $T=149360 121920 1 0 $X=149070 $Y=117710
X1642 450 443 384 1155 412 1 2 AOI31D0BWP7T $T=213760 114080 0 180 $X=210110 $Y=109870
X1643 913 1 36 12 2 38 ND3D0BWP7T $T=28400 121920 0 0 $X=28110 $Y=121685
X1644 326 1 389 357 2 1156 ND3D0BWP7T $T=195280 145440 0 0 $X=194990 $Y=145205
X1645 37 1 2 963 110 965 99 NR4D0BWP7T $T=56960 114080 0 0 $X=56670 $Y=113845
X1646 131 1 2 138 121 975 73 NR4D0BWP7T $T=67600 114080 1 180 $X=63950 $Y=113845
X1647 144 1 2 961 131 983 155 NR4D0BWP7T $T=69840 114080 1 0 $X=69550 $Y=109870
X1648 295 1 2 1033 289 1078 285 NR4D0BWP7T $T=135920 106240 1 180 $X=132270 $Y=106005
X1649 320 1 2 1055 334 1118 333 NR4D0BWP7T $T=153280 106240 1 180 $X=149630 $Y=106005
X1650 1160 1 2 426 425 1153 422 NR4D0BWP7T $T=197520 106240 1 180 $X=193870 $Y=106005
X1651 4 25 2 29 1 NR2D2BWP7T $T=23920 161120 0 0 $X=23630 $Y=160885
X1652 949 86 2 92 1 NR2D2BWP7T $T=51360 168960 1 0 $X=51070 $Y=164750
X1653 95 102 2 86 1 NR2D2BWP7T $T=58080 145440 1 180 $X=53870 $Y=145205
X1654 95 923 2 177 1 NR2D2BWP7T $T=85520 161120 0 0 $X=85230 $Y=160885
X1655 248 249 216 253 2 1 1044 AN4D1BWP7T $T=110720 137600 1 0 $X=110430 $Y=133390
X1656 1107 1 2 1108 BUFFD0BWP7T $T=151600 137600 0 180 $X=149070 $Y=133390
X1657 928 23 40 927 935 2 1 AOI31D1BWP7T $T=38480 121920 0 0 $X=38190 $Y=121685
X1658 965 969 979 142 982 2 1 AOI31D1BWP7T $T=67040 121920 0 0 $X=66750 $Y=121685
X1659 95 159 981 57 973 2 1 AOI31D1BWP7T $T=81600 145440 0 0 $X=81310 $Y=145205
X1660 1024 266 1053 1058 1060 2 1 AOI31D1BWP7T $T=122480 129760 0 0 $X=122190 $Y=129525
X1661 217 48 271 1011 25 2 1 AOI31D1BWP7T $T=123040 168960 1 0 $X=122750 $Y=164750
X1662 1177 1175 1148 445 412 2 1 AOI31D1BWP7T $T=218800 106240 1 180 $X=214590 $Y=106005
X1663 38 1 65 940 943 945 2 ND4D0BWP7T $T=44640 121920 0 0 $X=44350 $Y=121685
X1664 81 1 42 52 87 956 2 ND4D0BWP7T $T=50240 106240 0 0 $X=49950 $Y=106005
X1665 954 1 942 100 91 960 2 ND4D0BWP7T $T=54720 114080 1 0 $X=54430 $Y=109870
X1666 97 1 56 969 112 972 2 ND4D0BWP7T $T=60880 129760 1 0 $X=60590 $Y=125550
X1667 97 1 80 957 132 134 2 ND4D0BWP7T $T=62000 106240 0 0 $X=61710 $Y=106005
X1668 136 1 920 139 91 988 2 ND4D0BWP7T $T=65360 106240 0 0 $X=65070 $Y=106005
X1669 218 1 216 214 211 1021 2 ND4D0BWP7T $T=103440 114080 1 180 $X=99790 $Y=113845
X1670 219 1 1027 223 226 1028 2 ND4D0BWP7T $T=102880 121920 0 0 $X=102590 $Y=121685
X1671 231 1 236 1027 202 1034 2 ND4D0BWP7T $T=106240 121920 1 0 $X=105950 $Y=117710
X1672 216 1 236 214 1029 1040 2 ND4D0BWP7T $T=108480 129760 1 0 $X=108190 $Y=125550
X1673 247 1 240 250 251 1046 2 ND4D0BWP7T $T=110720 121920 1 0 $X=110430 $Y=117710
X1674 213 1 307 304 226 1090 2 ND4D0BWP7T $T=138720 106240 0 0 $X=138430 $Y=106005
X1675 444 1 442 441 439 1158 2 ND4D0BWP7T $T=213760 106240 1 180 $X=210110 $Y=106005
X1676 915 267 938 2 1 NR2D1P5BWP7T $T=121920 161120 0 0 $X=121630 $Y=160885
X1677 1019 1042 299 2 1 NR2D1P5BWP7T $T=134800 153280 0 0 $X=134510 $Y=153045
X1678 341 1137 399 2 1 NR2D1P5BWP7T $T=181840 153280 0 0 $X=181550 $Y=153045
X1679 436 440 430 2 1 NR2D1P5BWP7T $T=209280 121920 1 0 $X=208990 $Y=117710
X1680 499 1290 1321 2 1 NR2D1P5BWP7T $T=356000 114080 1 180 $X=351790 $Y=113845
X1681 54 2 932 64 68 942 1 INR4D0BWP7T $T=42960 114080 1 0 $X=42670 $Y=109870
X1682 5 2 71 947 941 943 1 INR4D0BWP7T $T=51360 121920 0 180 $X=46590 $Y=117710
X1683 82 2 85 935 922 958 1 INR4D0BWP7T $T=49680 114080 0 0 $X=49390 $Y=113845
X1684 228 1 1025 257 1043 2 NR3D1BWP7T $T=115200 114080 0 180 $X=110430 $Y=109870
X1685 278 1 283 1040 1068 2 NR3D1BWP7T $T=126960 129760 1 0 $X=126670 $Y=125550
X1686 208 1 202 200 1014 187 2 IND4D0BWP7T $T=100080 114080 1 180 $X=95870 $Y=113845
X1687 1038 1 1052 1081 1080 292 2 IND4D0BWP7T $T=138720 129760 0 180 $X=134510 $Y=125550
X1688 290 1 1109 346 1121 1122 2 IND4D0BWP7T $T=153280 114080 0 0 $X=152990 $Y=113845
X1689 208 1 236 243 1033 1037 2 IND4D1BWP7T $T=106240 114080 1 0 $X=105950 $Y=109870
X1690 946 2 79 93 949 1 103 NR4D3BWP7T $T=45200 153280 0 0 $X=44910 $Y=153045
X1691 1129 2 1136 1137 396 1 407 NR4D3BWP7T $T=175680 121920 1 0 $X=175390 $Y=117710
X1692 114 117 101 940 96 1 2 INR4D1BWP7T $T=60880 121920 0 180 $X=53870 $Y=117710
X1693 204 1016 210 1020 220 1 2 INR4D1BWP7T $T=97280 129760 1 0 $X=96990 $Y=125550
X1694 3 2 15 1 8 NR2XD1BWP7T $T=22240 145440 0 0 $X=21950 $Y=145205
X1695 13 2 35 1 44 NR2XD1BWP7T $T=41840 129760 0 0 $X=41550 $Y=129525
X1696 19 2 75 1 939 NR2XD1BWP7T $T=46320 129760 0 0 $X=46030 $Y=129525
X1697 952 2 115 1 973 NR2XD1BWP7T $T=62560 137600 0 0 $X=62270 $Y=137365
X1698 930 2 949 1 985 NR2XD1BWP7T $T=67040 153280 1 0 $X=66750 $Y=149070
X1699 4 2 152 1 985 NR2XD1BWP7T $T=69280 161120 0 0 $X=68990 $Y=160885
X1700 915 2 166 1 102 NR2XD1BWP7T $T=82160 161120 1 0 $X=81870 $Y=156910
X1701 915 2 167 1 4 NR2XD1BWP7T $T=82160 168960 1 0 $X=81870 $Y=164750
X1702 1001 2 171 1 176 NR2XD1BWP7T $T=84400 137600 1 0 $X=84110 $Y=133390
X1703 182 2 180 1 923 NR2XD1BWP7T $T=91120 161120 0 180 $X=86910 $Y=156910
X1704 159 2 169 1 163 NR2XD1BWP7T $T=91680 145440 1 180 $X=87470 $Y=145205
X1705 930 2 192 1 182 NR2XD1BWP7T $T=95600 161120 0 180 $X=91390 $Y=156910
X1706 1015 2 194 1 189 NR2XD1BWP7T $T=96720 106240 1 180 $X=92510 $Y=106005
X1707 176 2 966 1 195 NR2XD1BWP7T $T=100080 137600 0 180 $X=95870 $Y=133390
X1708 971 2 143 1 1023 NR2XD1BWP7T $T=97840 145440 0 0 $X=97550 $Y=145205
X1709 1039 2 250 1 1016 NR2XD1BWP7T $T=115200 121920 1 180 $X=110990 $Y=121685
X1710 1072 2 308 1 238 NR2XD1BWP7T $T=142640 161120 1 180 $X=138430 $Y=160885
X1711 1105 2 1101 1 1117 NR2XD1BWP7T $T=156640 145440 0 180 $X=152430 $Y=141230
X1712 332 2 1054 1 1105 NR2XD1BWP7T $T=157200 145440 1 180 $X=152990 $Y=145205
X1713 578 1 1286 579 2 IND2D1BWP7T $T=320720 168960 0 180 $X=317630 $Y=164750
X1714 232 233 225 239 2 1 1035 OR4XD1BWP7T $T=105680 106240 0 0 $X=105390 $Y=106005
X1715 1115 1113 1053 1102 2 1 348 OR4XD1BWP7T $T=151600 129760 1 0 $X=151310 $Y=125550
X1716 375 352 415 416 421 1 2 AO211D2BWP7T $T=189680 161120 0 0 $X=189390 $Y=160885
X1717 82 1 953 16 2 939 951 OAI211D0BWP7T $T=54160 129760 1 180 $X=50510 $Y=129525
X1718 82 1 953 16 2 939 959 OAI211D0BWP7T $T=58080 129760 1 180 $X=54430 $Y=129525
X1719 82 1 953 16 2 939 964 OAI211D0BWP7T $T=56960 129760 1 0 $X=56670 $Y=125550
X1720 375 1 381 350 2 341 1131 OAI211D0BWP7T $T=176240 161120 0 180 $X=172590 $Y=156910
X1721 1171 1 1145 388 2 385 1179 OAI211D0BWP7T $T=216000 145440 0 0 $X=215710 $Y=145205
X1722 597 1 1291 484 2 1296 1292 OAI211D0BWP7T $T=333040 114080 0 0 $X=332750 $Y=113845
X1723 633 1 1323 1325 2 1195 1310 OAI211D0BWP7T $T=358240 161120 0 180 $X=354590 $Y=156910
X1724 366 1 365 357 1126 1119 2 OAI211D2BWP7T $T=171760 145440 0 180 $X=165310 $Y=141230
X1725 433 1 432 365 1165 350 2 OAI211D2BWP7T $T=206480 161120 0 0 $X=206190 $Y=160885
X1726 1154 1 432 431 1168 399 2 OAI211D2BWP7T $T=207600 153280 0 0 $X=207310 $Y=153045
X1727 1171 1 1145 385 1187 388 2 OAI211D2BWP7T $T=217680 145440 1 0 $X=217390 $Y=141230
X1728 1222 1 1284 1195 570 576 2 OAI211D2BWP7T $T=315120 153280 0 180 $X=308670 $Y=149070
X1729 388 1 437 413 2 CKND2D3BWP7T $T=212080 129760 1 180 $X=206750 $Y=129525
X1730 22 23 932 47 1 2 929 AO211D0BWP7T $T=37920 114080 0 0 $X=37630 $Y=113845
X1731 1036 241 145 230 1 2 227 AO211D0BWP7T $T=109600 161120 1 180 $X=105390 $Y=160885
X1732 264 1054 1056 1057 1 2 1061 AO211D0BWP7T $T=123040 137600 0 0 $X=122750 $Y=137365
X1733 429 431 1161 1159 1 2 1163 AO211D0BWP7T $T=205920 153280 1 0 $X=205630 $Y=149070
X1734 466 1219 1199 1260 1 2 1262 AO211D0BWP7T $T=292160 153280 1 0 $X=291870 $Y=149070
X1735 979 2 179 994 966 1000 1 AOI211D2BWP7T $T=90560 129760 0 180 $X=84110 $Y=125550
X1736 917 2 11 13 1 NR2D3BWP7T $T=28400 145440 0 180 $X=23070 $Y=141230
X1737 915 2 32 923 1 NR2D3BWP7T $T=23360 153280 0 0 $X=23070 $Y=153045
X1738 962 2 83 971 1 NR2D3BWP7T $T=59200 145440 1 0 $X=58910 $Y=141230
X1739 952 2 93 102 1 NR2D3BWP7T $T=67040 153280 0 180 $X=61710 $Y=149070
X1740 930 2 145 984 1 NR2D3BWP7T $T=65360 145440 0 0 $X=65070 $Y=145205
X1741 923 2 160 57 1 NR2D3BWP7T $T=84960 161120 1 180 $X=79630 $Y=160885
X1742 95 2 191 1011 1 NR2D3BWP7T $T=89440 161120 0 0 $X=89150 $Y=160885
X1743 95 2 230 4 1 NR2D3BWP7T $T=112960 168960 0 180 $X=107630 $Y=164750
X1744 1051 2 272 238 1 NR2D3BWP7T $T=129200 145440 1 180 $X=123870 $Y=145205
X1745 1019 2 229 273 1 NR2D3BWP7T $T=131440 153280 1 180 $X=126110 $Y=153045
X1746 336 2 339 345 1 NR2D3BWP7T $T=149920 153280 0 0 $X=149630 $Y=153045
X1747 341 2 344 337 1 NR2D3BWP7T $T=152160 168960 1 0 $X=151870 $Y=164750
X1748 350 2 429 388 1 NR2D3BWP7T $T=210960 137600 0 0 $X=210670 $Y=137365
X1749 242 1023 1 2 107 AN2D1BWP7T $T=108480 153280 0 0 $X=108190 $Y=153045
X1750 429 1156 1 2 1173 AN2D1BWP7T $T=214320 129760 0 0 $X=214030 $Y=129525
X1751 916 19 15 1 2 ND2D2BWP7T $T=30080 129760 1 180 $X=25870 $Y=129525
X1752 35 28 928 1 2 ND2D2BWP7T $T=41840 129760 1 180 $X=37630 $Y=129525
X1753 933 41 49 1 2 ND2D2BWP7T $T=41840 137600 1 180 $X=37630 $Y=137365
X1754 107 95 971 1 2 ND2D2BWP7T $T=69280 145440 0 180 $X=65070 $Y=141230
X1755 242 57 143 1 2 ND2D2BWP7T $T=110720 153280 0 180 $X=106510 $Y=149070
X1756 238 923 1042 1 2 ND2D2BWP7T $T=113520 145440 0 180 $X=109310 $Y=141230
X1757 242 915 1041 1 2 ND2D2BWP7T $T=114640 153280 0 180 $X=110430 $Y=149070
X1758 1041 182 221 1 2 ND2D2BWP7T $T=110720 161120 1 0 $X=110430 $Y=156910
X1759 273 102 1077 1 2 ND2D2BWP7T $T=134800 161120 0 180 $X=130590 $Y=156910
X1760 308 48 299 1 2 ND2D2BWP7T $T=138720 168960 1 0 $X=138430 $Y=164750
X1761 368 328 341 1 2 ND2D2BWP7T $T=171200 153280 1 180 $X=166990 $Y=153045
X1762 388 387 362 1 2 ND2D2BWP7T $T=176240 168960 1 0 $X=175950 $Y=164750
X1763 436 412 430 1 2 ND2D2BWP7T $T=217680 114080 1 180 $X=213470 $Y=113845
X1764 446 531 1184 1 2 ND2D2BWP7T $T=279280 153280 0 0 $X=278990 $Y=153045
X1765 561 2 1272 1258 542 1 571 1274 AOI221D1BWP7T $T=305600 153280 0 0 $X=305310 $Y=153045
X1766 113 1 2 73 99 120 NR3D0BWP7T $T=59200 106240 0 0 $X=58910 $Y=106005
X1767 115 1 2 949 119 118 NR3D0BWP7T $T=59200 168960 1 0 $X=58910 $Y=164750
X1768 1005 1 2 166 119 172 NR3D0BWP7T $T=88880 168960 0 180 $X=85790 $Y=164750
X1769 261 1 2 262 1026 1052 NR3D0BWP7T $T=121920 121920 0 0 $X=121630 $Y=121685
X1770 1099 1097 1 1073 1098 2 AOI21D1BWP7T $T=144320 137600 1 180 $X=140670 $Y=137365
X1771 1099 1080 1 1093 317 2 AOI21D1BWP7T $T=144880 145440 1 180 $X=141230 $Y=145205
X1772 353 368 1 337 1139 2 AOI21D1BWP7T $T=184080 161120 0 0 $X=183790 $Y=160885
X1773 477 586 1 1289 1284 2 AOI21D1BWP7T $T=317920 153280 1 0 $X=317630 $Y=149070
X1774 621 620 1 1303 1307 2 AOI21D1BWP7T $T=347040 114080 0 180 $X=343390 $Y=109870
X1775 8 3 18 916 2 1 ND3D2BWP7T $T=21120 129760 0 0 $X=20830 $Y=129525
X1776 8 12 62 3 2 1 ND3D2BWP7T $T=42960 153280 1 0 $X=42670 $Y=149070
X1777 258 2 1025 1037 1 NR2D0BWP7T $T=114640 106240 1 180 $X=112110 $Y=106005
X1778 112 1 961 14 913 916 2 OAI31D2BWP7T $T=59200 137600 1 180 $X=52190 $Y=137365
X1779 966 1 976 972 918 126 2 OAI31D2BWP7T $T=69280 129760 1 180 $X=62270 $Y=129525
X1780 1101 1 1104 373 1123 364 2 OAI31D2BWP7T $T=166160 121920 1 0 $X=165870 $Y=117710
X1781 1029 1 248 1043 2 255 ND3D1BWP7T $T=111840 129760 0 0 $X=111550 $Y=129525
X1782 1201 2 484 1198 1 1196 478 AOI211D1BWP7T $T=237840 145440 0 180 $X=234190 $Y=141230
X1783 483 2 484 488 1 491 493 AOI211D1BWP7T $T=235600 168960 1 0 $X=235310 $Y=164750
X1784 518 2 1228 519 1 1221 482 AOI211D1BWP7T $T=267520 106240 0 0 $X=267230 $Y=106005
X1785 1336 2 1290 1330 1 1331 466 AOI211D1BWP7T $T=367200 114080 1 180 $X=363550 $Y=113845
X1786 1340 2 659 1338 1 1323 482 AOI211D1BWP7T $T=378960 153280 0 180 $X=375310 $Y=149070
X1787 1347 2 1290 1343 1 1342 466 AOI211D1BWP7T $T=382320 121920 0 180 $X=378670 $Y=117710
X1788 1376 2 682 1375 1 1372 466 AOI211D1BWP7T $T=407520 121920 0 180 $X=403870 $Y=117710
X1789 711 743 714 749 736 1 2 758 AO221D0BWP7T $T=436080 129760 0 0 $X=435790 $Y=129525
X1790 712 744 717 1386 736 1 2 1387 AO221D0BWP7T $T=440560 114080 1 0 $X=440270 $Y=109870
X1813 374 1216 382 1207 2 1 501 DFCND1BWP7T $T=263600 153280 1 180 $X=250430 $Y=153045
X1814 374 1316 605 1326 2 1 643 DFCND1BWP7T $T=349280 145440 0 0 $X=348990 $Y=145205
X1815 475 468 464 1 2 XNR2D2BWP7T $T=233920 145440 1 180 $X=226910 $Y=145205
X1816 987 1 2 170 956 1004 105 AOI211XD0BWP7T $T=84960 114080 1 0 $X=84670 $Y=109870
X1817 152 1 2 209 1019 1018 124 AOI211XD0BWP7T $T=101760 168960 0 180 $X=98110 $Y=164750
X1818 198 1 2 145 1030 235 237 AOI211XD0BWP7T $T=104560 168960 1 0 $X=104270 $Y=164750
X1819 1096 1 2 1089 1065 1092 1062 AOI211XD0BWP7T $T=142640 114080 1 180 $X=138990 $Y=113845
X1820 404 1 2 1140 402 1142 378 AOI211XD0BWP7T $T=187440 114080 0 180 $X=183790 $Y=109870
X1821 1196 1 2 1199 1198 479 466 AOI211XD0BWP7T $T=237840 153280 0 180 $X=234190 $Y=149070
X1822 1247 1 2 1253 540 1245 482 AOI211XD0BWP7T $T=290480 106240 0 0 $X=290190 $Y=106005
X1823 1324 1 2 1322 1314 1308 482 AOI211XD0BWP7T $T=358240 145440 0 180 $X=354590 $Y=141230
X1824 374 1217 382 504 502 1 2 DFCND2BWP7T $T=264720 161120 1 180 $X=249870 $Y=160885
X1825 374 1212 382 1214 1229 1 2 DFCND2BWP7T $T=252960 129760 1 0 $X=252670 $Y=125550
X1826 374 1320 525 1313 1311 1 2 DFCND2BWP7T $T=362160 129760 0 180 $X=347310 $Y=125550
X1827 374 1368 525 667 1351 1 2 DFCND2BWP7T $T=404160 129760 0 180 $X=389310 $Y=125550
X1828 50 1 61 938 57 2 OAI21D2BWP7T $T=40720 168960 1 0 $X=40430 $Y=164750
X1829 188 1 197 984 1011 2 OAI21D2BWP7T $T=91680 168960 1 0 $X=91390 $Y=164750
X1830 399 389 1 351 2 1159 381 OAI22D1BWP7T $T=194160 161120 1 0 $X=193870 $Y=156910
X1831 336 326 1 365 2 428 350 OAI22D1BWP7T $T=194720 168960 1 0 $X=194430 $Y=164750
X1832 326 417 1 435 2 1161 388 OAI22D1BWP7T $T=205920 168960 1 0 $X=205630 $Y=164750
X1833 603 545 1 543 2 1289 1300 OAI22D1BWP7T $T=335840 137600 1 0 $X=335550 $Y=133390
X1834 1004 1 2 1007 DEL1BWP7T $T=95600 114080 1 180 $X=89710 $Y=113845
X1835 549 560 550 1270 561 1 2 569 AO221D1BWP7T $T=303920 137600 1 0 $X=303630 $Y=133390
X1836 541 572 1251 1278 578 1 2 1280 AO221D1BWP7T $T=308960 114080 1 0 $X=308670 $Y=109870
X1837 596 1293 599 1297 561 1 2 607 AO221D1BWP7T $T=333040 137600 0 0 $X=332750 $Y=137365
X1838 1295 530 1191 1299 578 1 2 614 AO221D1BWP7T $T=335280 129760 1 0 $X=334990 $Y=125550
X1839 595 600 598 1294 578 1 2 615 AO221D1BWP7T $T=336400 114080 1 0 $X=336110 $Y=109870
X1840 594 609 1226 1301 578 1 2 1302 AO221D1BWP7T $T=336960 161120 0 0 $X=336670 $Y=160885
X1841 680 715 678 1377 578 1 2 720 AO221D1BWP7T $T=417600 137600 0 0 $X=417310 $Y=137365
X1842 676 708 1333 1382 578 1 2 1384 AO221D1BWP7T $T=421520 153280 0 0 $X=421230 $Y=153045
X1843 721 658 1383 1380 578 1 2 734 AO221D1BWP7T $T=422640 145440 1 0 $X=422350 $Y=141230
X1844 374 1205 382 512 2 1 1211 DFCND0BWP7T $T=247920 137600 1 0 $X=247630 $Y=133390
X1845 374 1206 382 1204 2 1 513 DFCND0BWP7T $T=249040 121920 0 0 $X=248750 $Y=121685
X1846 374 1210 382 1218 2 1 1224 DFCND0BWP7T $T=252400 129760 0 0 $X=252110 $Y=129525
X1847 374 515 382 520 2 1 1237 DFCND0BWP7T $T=259680 168960 1 0 $X=259390 $Y=164750
X1848 374 1231 382 1238 2 1 1241 DFCND0BWP7T $T=266960 121920 0 0 $X=266670 $Y=121685
X1849 374 1232 525 1234 2 1 1190 DFCND0BWP7T $T=282080 161120 0 180 $X=268910 $Y=156910
X1850 374 1215 525 1240 2 1 534 DFCND0BWP7T $T=269760 114080 1 0 $X=269470 $Y=109870
X1851 374 1233 525 1239 2 1 1389 DFCND0BWP7T $T=269760 145440 1 0 $X=269470 $Y=141230
X1852 374 1244 525 1235 2 1 1225 DFCND0BWP7T $T=283200 137600 0 180 $X=270030 $Y=133390
X1853 374 1257 525 1252 2 1 1265 DFCND0BWP7T $T=291040 121920 0 0 $X=290750 $Y=121685
X1854 374 1256 525 548 2 1 1269 DFCND0BWP7T $T=292160 114080 0 0 $X=291870 $Y=113845
X1855 374 1267 525 1275 2 1 1276 DFCND0BWP7T $T=297760 106240 0 0 $X=297470 $Y=106005
X1856 374 1315 605 1327 2 1 1390 DFCND0BWP7T $T=349280 153280 0 0 $X=348990 $Y=153045
X1857 374 1328 525 1318 2 1 1309 DFCND0BWP7T $T=363840 121920 1 180 $X=350670 $Y=121685
X1858 374 1360 525 665 2 1 1352 DFCND0BWP7T $T=399120 106240 1 180 $X=385950 $Y=106005
X1859 374 1362 605 1356 2 1 1354 DFCND0BWP7T $T=402480 145440 0 180 $X=389310 $Y=141230
X1860 374 1357 605 1355 2 1 1344 DFCND0BWP7T $T=402480 161120 0 180 $X=389310 $Y=156910
X1861 1191 506 474 507 480 510 2 1213 1 OA222D0BWP7T $T=252400 121920 1 0 $X=252110 $Y=117710
X1862 516 506 388 1218 503 512 2 1208 1 OA222D0BWP7T $T=264160 137600 1 180 $X=257710 $Y=137365
X1863 524 506 388 1235 503 1218 2 1227 1 OA222D0BWP7T $T=275360 137600 1 180 $X=268910 $Y=137365
X1864 1242 506 388 523 503 1238 2 1236 1 OA222D0BWP7T $T=277600 129760 1 180 $X=271150 $Y=129525
X1865 1258 506 526 520 503 1252 2 1250 1 OA222D0BWP7T $T=296080 145440 1 180 $X=289630 $Y=145205
X1866 1254 555 526 1238 503 548 2 1259 1 OA222D0BWP7T $T=302800 114080 0 180 $X=296350 $Y=109870
X1867 651 640 526 644 503 632 2 639 1 OA222D0BWP7T $T=366080 168960 0 180 $X=359630 $Y=164750
X1868 694 640 526 1355 503 681 2 679 1 OA222D0BWP7T $T=397440 168960 0 180 $X=390990 $Y=164750
X1869 701 640 526 661 503 693 2 1363 1 OA222D0BWP7T $T=404160 153280 1 180 $X=397710 $Y=153045
X1870 924 2 37 1 920 914 22 AOI211XD1BWP7T $T=31200 114080 1 180 $X=24190 $Y=113845
X1871 93 2 166 1 183 163 175 AOI211XD1BWP7T $T=82720 153280 0 0 $X=82430 $Y=153045
X1872 339 2 405 1 1151 359 414 AOI211XD1BWP7T $T=186320 168960 1 0 $X=186030 $Y=164750
X1873 927 13 1 2 INVD2P5BWP7T $T=31200 145440 0 180 $X=28110 $Y=141230
X1874 602 606 1 2 INVD2P5BWP7T $T=335280 161120 1 0 $X=334990 $Y=156910
X1875 1286 612 1 2 INVD2P5BWP7T $T=337520 153280 0 0 $X=337230 $Y=153045
X1876 1388 787 1 2 INVD2P5BWP7T $T=464080 153280 1 0 $X=463790 $Y=149070
X1877 783 792 1 2 INVD2P5BWP7T $T=466320 121920 1 0 $X=466030 $Y=117710
X1878 790 795 1 2 INVD2P5BWP7T $T=466320 161120 0 0 $X=466030 $Y=160885
X1879 799 801 1 2 INVD2P5BWP7T $T=473040 161120 1 180 $X=469950 $Y=160885
X1880 381 388 1 2 INVD6BWP7T $T=213200 137600 0 180 $X=207870 $Y=133390
X1881 506 514 1 474 500 503 508 2 1206 OAI222D2BWP7T $T=261360 114080 0 180 $X=250990 $Y=109870
X1882 506 511 1 474 504 503 500 2 1217 OAI222D2BWP7T $T=263600 161120 0 180 $X=253230 $Y=156910
X1883 506 1226 1 474 1207 503 1214 2 1216 OAI222D2BWP7T $T=265280 153280 0 180 $X=254910 $Y=149070
X1884 506 1243 1 388 1234 503 521 2 1232 OAI222D2BWP7T $T=279840 161120 1 180 $X=269470 $Y=160885
X1885 506 1251 1 474 1214 503 522 2 1212 OAI222D2BWP7T $T=280400 114080 1 180 $X=270030 $Y=113845
X1886 506 533 1 526 452 503 1234 2 1233 OAI222D2BWP7T $T=280400 153280 0 180 $X=270030 $Y=149070
X1887 506 552 1 526 1235 503 1252 2 1244 OAI222D2BWP7T $T=300560 137600 1 180 $X=290190 $Y=137365
X1888 640 648 1 526 630 503 1313 2 1315 OAI222D2BWP7T $T=362160 161120 1 180 $X=351790 $Y=160885
X1889 640 1333 1 526 1326 503 632 2 1316 OAI222D2BWP7T $T=363840 153280 0 180 $X=353470 $Y=149070
X1890 640 647 1 526 1313 503 635 2 1320 OAI222D2BWP7T $T=364960 129760 1 180 $X=354590 $Y=129525
X1891 640 650 1 526 626 503 637 2 1328 OAI222D2BWP7T $T=366080 137600 0 180 $X=355710 $Y=133390
X1892 555 700 1 526 667 503 686 2 1368 OAI222D2BWP7T $T=403600 114080 1 180 $X=393230 $Y=113845
X1893 640 1373 1 526 1355 503 690 2 1357 OAI222D2BWP7T $T=403600 153280 0 180 $X=393230 $Y=149070
X1894 429 1 2 336 INVD5BWP7T $T=211520 145440 0 180 $X=206750 $Y=141230
X1895 927 2 1 66 60 NR2D2P5BWP7T $T=50240 137600 1 180 $X=44910 $Y=137365
X1896 238 229 175 2 1 CKAN2D2BWP7T $T=107920 145440 1 180 $X=103710 $Y=145205
X1897 163 992 1 2 153 CKAN2D1BWP7T $T=82720 153280 1 180 $X=79630 $Y=153045
X1898 1112 1059 1103 1088 2 1 340 AN4D0BWP7T $T=149360 121920 0 0 $X=149070 $Y=121685
X1899 950 2 70 936 77 1 NR3D2BWP7T $T=52480 161120 0 180 $X=42110 $Y=156910
X1900 19 14 5 1 2 OR2D2BWP7T $T=25040 121920 0 180 $X=20830 $Y=117710
X1901 12 16 6 1 2 OR2D2BWP7T $T=25600 106240 1 180 $X=21390 $Y=106005
X1902 8 9 7 1 2 OR2D2BWP7T $T=25600 121920 1 180 $X=21390 $Y=121685
X1903 242 270 25 1 2 OR2D2BWP7T $T=124160 161120 1 0 $X=123870 $Y=156910
X1904 1185 417 461 1 2 OR2D2BWP7T $T=223280 137600 0 0 $X=222990 $Y=137365
X1905 49 66 44 1 2 ND2D1P5BWP7T $T=46320 145440 1 0 $X=46030 $Y=141230
X1906 18 23 1 2 INVD1P5BWP7T $T=23920 129760 1 0 $X=23630 $Y=125550
X1907 86 2 79 107 1 108 20 AOI211XD2BWP7T $T=49120 153280 1 0 $X=48830 $Y=149070
X1908 1108 2 1111 1114 1 343 1101 AOI211XD2BWP7T $T=144320 137600 0 0 $X=144030 $Y=137365
X1909 1282 2 1290 582 1 590 466 AOI211XD2BWP7T $T=324640 129760 0 180 $X=311470 $Y=125550
X1910 1307 2 631 620 1 623 466 AOI211XD2BWP7T $T=354320 106240 1 180 $X=341150 $Y=106005
X1911 689 2 682 1366 1 699 466 AOI211XD2BWP7T $T=393520 114080 1 0 $X=393230 $Y=109870
X1912 984 2 1 119 923 NR2XD2BWP7T $T=83280 153280 1 0 $X=82990 $Y=149070
X1913 102 2 1 199 984 NR2XD2BWP7T $T=101200 153280 1 180 $X=94190 $Y=153045
X1914 387 2 1 1138 328 NR2XD2BWP7T $T=179040 161120 1 0 $X=178750 $Y=156910
X1915 1 2 ICV_23 $T=27280 121920 1 0 $X=26990 $Y=117710
X1916 1 2 ICV_23 $T=69280 145440 1 0 $X=68990 $Y=141230
X1917 1 2 ICV_23 $T=153280 106240 0 0 $X=152990 $Y=106005
X1918 1 2 ICV_23 $T=193600 121920 0 0 $X=193310 $Y=121685
X1919 1 2 ICV_23 $T=263600 153280 0 0 $X=263310 $Y=153045
X1920 1 2 ICV_23 $T=277600 129760 0 0 $X=277310 $Y=129525
X1921 1 2 ICV_23 $T=308960 145440 0 0 $X=308670 $Y=145205
X1922 1 2 ICV_23 $T=321280 161120 0 0 $X=320990 $Y=160885
X1923 1 2 ICV_23 $T=342560 161120 0 0 $X=342270 $Y=160885
X1924 1 2 ICV_23 $T=371120 114080 1 0 $X=370830 $Y=109870
X1925 1 2 ICV_23 $T=403600 114080 0 0 $X=403310 $Y=113845
X1926 1 2 ICV_23 $T=413120 153280 1 0 $X=412830 $Y=149070
X1927 1 2 ICV_23 $T=445600 114080 1 0 $X=445310 $Y=109870
X1928 1 2 ICV_23 $T=445600 114080 0 0 $X=445310 $Y=113845
X1929 1 2 ICV_23 $T=445600 129760 1 0 $X=445310 $Y=125550
X1930 1 2 ICV_23 $T=447280 153280 1 0 $X=446990 $Y=149070
X1931 1 2 ICV_23 $T=455120 153280 1 0 $X=454830 $Y=149070
X1932 1 2 ICV_23 $T=465760 129760 1 0 $X=465470 $Y=125550
X1933 476 526 1 2 INVD8BWP7T $T=293840 129760 0 0 $X=293550 $Y=129525
X1934 931 12 8 53 1 2 AN3D2BWP7T $T=39600 145440 0 0 $X=39310 $Y=145205
X1935 44 49 927 14 2 1 OR3D2BWP7T $T=50800 145440 1 0 $X=50510 $Y=141230
X1936 974 994 920 995 991 994 2 1 AOI32D1BWP7T $T=79920 129760 1 0 $X=79630 $Y=125550
X1937 977 1007 150 1009 133 1004 2 1 AOI32D1BWP7T $T=92800 121920 0 180 $X=88030 $Y=117710
X1938 357 359 353 1124 351 350 2 1 AOI32D1BWP7T $T=168400 161120 0 180 $X=163630 $Y=156910
X1939 345 350 328 1127 359 385 2 1 AOI32D1BWP7T $T=172880 153280 0 0 $X=172590 $Y=153045
X1958 537 564 1243 492 561 575 1 2 AO221D2BWP7T $T=305600 161120 0 0 $X=305310 $Y=160885
X1959 683 727 688 733 578 735 1 2 AO221D2BWP7T $T=425440 168960 1 0 $X=425150 $Y=164750
X1960 336 1 326 1130 350 365 2 OAI22D2BWP7T $T=165600 145440 0 0 $X=165310 $Y=145205
X1961 1248 1 545 536 539 543 2 OAI22D2BWP7T $T=296640 168960 0 180 $X=289630 $Y=164750
X1962 1288 1 545 1282 1285 543 2 OAI22D2BWP7T $T=322960 129760 1 180 $X=315950 $Y=129525
X1963 1066 1064 1056 1060 274 2 1 OAI22D0BWP7T $T=130320 137600 0 180 $X=126670 $Y=133390
X1964 1094 325 1107 1060 1095 2 1 OAI22D0BWP7T $T=149360 137600 0 180 $X=145710 $Y=133390
X1965 1094 329 1096 1066 319 2 1 OAI22D0BWP7T $T=150480 114080 1 180 $X=146830 $Y=113845
X1966 545 1263 1260 543 1264 2 1 OAI22D0BWP7T $T=302240 153280 1 180 $X=298590 $Y=153045
X1967 545 1283 1281 461 1277 2 1 OAI22D0BWP7T $T=317920 137600 1 180 $X=314270 $Y=137365
X1968 921 21 1 2 BUFFD4BWP7T $T=28960 153280 0 180 $X=23630 $Y=149070
X1969 1141 350 1 2 BUFFD4BWP7T $T=189680 137600 0 0 $X=189390 $Y=137365
X1970 1139 446 1 2 BUFFD4BWP7T $T=212640 161120 0 0 $X=212350 $Y=160885
X1971 1181 381 1 2 BUFFD4BWP7T $T=221040 129760 0 180 $X=215710 $Y=125550
X1972 1186 474 1 2 BUFFD4BWP7T $T=228320 114080 0 0 $X=228030 $Y=113845
X1973 978 986 998 165 1 1006 2 ND4D4BWP7T $T=81040 137600 0 0 $X=80750 $Y=137365
X1974 761 762 765 1 2 AN2D2BWP7T $T=443920 137600 1 0 $X=443630 $Y=133390
X1975 561 2 1254 1 669 NR2XD3BWP7T $T=384560 145440 0 180 $X=375870 $Y=141230
X1976 578 2 719 1 730 NR2XD3BWP7T $T=429920 161120 0 180 $X=421230 $Y=156910
X1977 578 2 705 1 731 NR2XD3BWP7T $T=430480 161120 1 180 $X=421790 $Y=160885
X1978 736 2 694 1 732 NR2XD3BWP7T $T=431040 137600 0 180 $X=422350 $Y=133390
X1979 736 2 1373 1 742 NR2XD3BWP7T $T=436640 121920 1 180 $X=427950 $Y=121685
X1980 578 2 745 1 767 NR2XD3BWP7T $T=445600 161120 0 180 $X=436910 $Y=156910
X1981 578 2 752 1 763 NR2XD3BWP7T $T=446720 168960 0 180 $X=438030 $Y=164750
X1982 355 360 369 382 353 341 1 2 EDFCND2BWP7T $T=165600 161120 0 0 $X=165310 $Y=160885
X1983 355 352 374 382 359 1141 1 2 EDFCND2BWP7T $T=168400 137600 0 0 $X=168110 $Y=137365
X1984 355 367 369 382 368 375 1 2 EDFCND2BWP7T $T=168400 153280 1 0 $X=168110 $Y=149070
X1985 1106 2 1083 1087 1076 294 1 NR4D4BWP7T $T=152160 153280 0 180 $X=130590 $Y=149070
X1986 1125 2 376 1134 398 395 1 NR4D4BWP7T $T=166160 114080 0 0 $X=165870 $Y=113845
X1987 1126 2 380 1133 1138 400 1 NR4D4BWP7T $T=168400 129760 1 0 $X=168110 $Y=125550
X1988 1132 2 1135 1143 413 1144 1 NR4D4BWP7T $T=172320 121920 0 0 $X=172030 $Y=121685
X1989 1128 2 1130 339 1138 411 1 NR4D4BWP7T $T=172880 137600 1 0 $X=172590 $Y=133390
X1990 327 1 1086 2 1097 OR2D0BWP7T $T=146000 121920 1 180 $X=142910 $Y=121685
X1991 937 74 953 957 2 56 1 IINR4D1BWP7T $T=48000 121920 0 0 $X=47710 $Y=121685
X1992 561 2 1242 1 748 NR2D5BWP7T $T=443360 145440 0 180 $X=434670 $Y=141230
X1993 561 2 746 1 755 NR2D5BWP7T $T=445040 153280 1 180 $X=436350 $Y=153045
X1994 578 2 757 1 759 NR2D5BWP7T $T=447840 161120 1 180 $X=439150 $Y=160885
X1995 561 565 554 1 2 INR2XD4BWP7T $T=314000 145440 0 180 $X=300830 $Y=141230
X1996 736 740 729 1 2 INR2XD4BWP7T $T=440560 137600 1 180 $X=427390 $Y=137365
X1997 736 750 737 1 2 INR2XD4BWP7T $T=445600 114080 1 180 $X=432430 $Y=113845
X1998 736 751 706 1 2 INR2XD4BWP7T $T=445600 129760 0 180 $X=432430 $Y=125550
X1999 736 754 611 1 2 INR2XD4BWP7T $T=446160 106240 1 180 $X=432990 $Y=106005
X2000 561 753 741 1 2 INR2XD4BWP7T $T=446720 145440 1 180 $X=433550 $Y=145205
X2001 561 756 722 1 2 INR2XD4BWP7T $T=447280 153280 0 180 $X=434110 $Y=149070
X2002 736 760 747 1 2 INR2XD4BWP7T $T=450080 121920 1 180 $X=436910 $Y=121685
X2003 561 780 768 1 2 INR2XD4BWP7T $T=470800 145440 1 180 $X=457630 $Y=145205
X2004 561 784 770 1 2 INR2XD4BWP7T $T=471920 153280 1 180 $X=458750 $Y=153045
X2005 561 791 773 1 2 INR2XD4BWP7T $T=474160 129760 1 180 $X=460990 $Y=129525
X2006 561 789 772 1 2 INR2XD4BWP7T $T=474160 137600 1 180 $X=460990 $Y=137365
X2007 984 1 973 2 205 OR2D1BWP7T $T=96160 153280 1 0 $X=95870 $Y=149070
X2008 446 1 399 2 1178 OR2D1BWP7T $T=217120 161120 1 0 $X=216830 $Y=156910
X2009 709 1 578 2 1381 OR2D1BWP7T $T=417600 168960 1 0 $X=417310 $Y=164750
X2010 716 1 736 2 1385 OR2D1BWP7T $T=431600 114080 1 0 $X=431310 $Y=109870
X2011 1 2 ICV_31 $T=32320 153280 0 0 $X=32030 $Y=153045
X2012 1 2 ICV_31 $T=32320 161120 0 0 $X=32030 $Y=160885
X2013 1 2 ICV_31 $T=74320 168960 1 0 $X=74030 $Y=164750
X2014 1 2 ICV_31 $T=116320 114080 0 0 $X=116030 $Y=113845
X2015 1 2 ICV_31 $T=116320 121920 1 0 $X=116030 $Y=117710
X2016 1 2 ICV_31 $T=116320 129760 1 0 $X=116030 $Y=125550
X2017 1 2 ICV_31 $T=158320 137600 1 0 $X=158030 $Y=133390
X2018 1 2 ICV_31 $T=200320 161120 1 0 $X=200030 $Y=156910
X2019 1 2 ICV_31 $T=242320 114080 0 0 $X=242030 $Y=113845
X2020 1 2 ICV_31 $T=242320 121920 0 0 $X=242030 $Y=121685
X2021 1 2 ICV_31 $T=242320 145440 1 0 $X=242030 $Y=141230
X2022 1 2 ICV_31 $T=242320 153280 1 0 $X=242030 $Y=149070
X2023 1 2 ICV_31 $T=284320 121920 0 0 $X=284030 $Y=121685
X2024 1 2 ICV_31 $T=284320 129760 0 0 $X=284030 $Y=129525
X2025 1 2 ICV_31 $T=284320 161120 0 0 $X=284030 $Y=160885
X2026 1 2 ICV_31 $T=368320 121920 0 0 $X=368030 $Y=121685
X2027 1 2 ICV_31 $T=368320 153280 1 0 $X=368030 $Y=149070
X2028 1 2 ICV_31 $T=410320 114080 0 0 $X=410030 $Y=113845
X2029 1 2 ICV_31 $T=452320 114080 0 0 $X=452030 $Y=113845
X2030 1 2 ICV_31 $T=452320 121920 1 0 $X=452030 $Y=117710
X2031 1 2 ICV_31 $T=452320 137600 1 0 $X=452030 $Y=133390
X2032 1 2 ICV_31 $T=452320 161120 1 0 $X=452030 $Y=156910
X2033 1 2 ICV_31 $T=452320 161120 0 0 $X=452030 $Y=160885
X2034 1 2 ICV_31 $T=472480 129760 1 0 $X=472190 $Y=125550
X2035 341 1 326 337 2 ND2D3BWP7T $T=156080 161120 0 180 $X=150750 $Y=156910
X2036 350 1 399 381 2 ND2D3BWP7T $T=208720 145440 0 0 $X=208430 $Y=145205
.ENDS
***************************************
.SUBCKT ICV_33 1 2
** N=2 EP=2 IP=4 FDC=4
X1 1 2 ICV_3 $T=0 0 0 0 $X=-290 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_34 1 2
** N=2 EP=2 IP=4 FDC=8
X0 1 2 ICV_3 $T=0 0 0 0 $X=-290 $Y=-235
X1 1 2 ICV_8 $T=2800 0 0 0 $X=2510 $Y=-235
.ENDS
***************************************
.SUBCKT ICV_35 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480
+ 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500
+ 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520
+ 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540
+ 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560
+ 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580
+ 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600
+ 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620
+ 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640
+ 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660
+ 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680
+ 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700
+ 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720
+ 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740
+ 741 742 743 744 745 746 747 748 749
** N=1347 EP=749 IP=7212 FDC=9618
M0 1 921 925 1 N L=1.8e-07 W=5e-07 $X=95100 $Y=97400 $D=0
M1 196 925 1 1 N L=1.8e-07 W=5e-07 $X=95760 $Y=97080 $D=0
M2 1 914 196 1 N L=1.8e-07 W=5e-07 $X=96480 $Y=97080 $D=0
M3 1 972 986 1 N L=1.8e-07 W=5e-07 $X=137100 $Y=97400 $D=0
M4 986 289 1 1 N L=1.8e-07 W=5e-07 $X=138060 $Y=97400 $D=0
M5 1 1003 986 1 N L=1.8e-07 W=5e-07 $X=138880 $Y=97400 $D=0
M6 1003 288 1 1 N L=1.8e-07 W=4.2e-07 $X=139600 $Y=97480 $D=0
M7 2 921 925 2 P L=1.8e-07 W=6.85e-07 $X=95100 $Y=94825 $D=16
M8 1345 925 2 2 P L=1.8e-07 W=1.37e-06 $X=95880 $Y=94825 $D=16
M9 196 914 1345 2 P L=1.8e-07 W=1.37e-06 $X=96480 $Y=94825 $D=16
M10 1346 972 986 2 P L=1.8e-07 W=1.37e-06 $X=137100 $Y=94825 $D=16
M11 1347 289 1346 2 P L=1.8e-07 W=1.37e-06 $X=137940 $Y=94825 $D=16
M12 2 1003 1347 2 P L=1.8e-07 W=1.37e-06 $X=138780 $Y=94825 $D=16
M13 1003 288 2 2 P L=1.8e-07 W=4.2e-07 $X=139600 $Y=95510 $D=16
X206 817 1 2 38 CKBD1BWP7T $T=27840 67040 0 0 $X=27550 $Y=66805
X207 981 1 2 952 CKBD1BWP7T $T=129760 82720 1 180 $X=127230 $Y=82485
X208 1230 1 2 1148 CKBD1BWP7T $T=278720 90560 0 180 $X=276190 $Y=86350
X209 570 1 2 1262 CKBD1BWP7T $T=331920 90560 1 0 $X=331630 $Y=86350
X210 1270 1 2 593 CKBD1BWP7T $T=353200 106240 0 180 $X=350670 $Y=102030
X211 603 1 2 634 CKBD1BWP7T $T=390720 90560 1 180 $X=388190 $Y=90325
X212 638 1 2 641 CKBD1BWP7T $T=392400 106240 1 0 $X=392110 $Y=102030
X213 808 1 2 823 INVD0BWP7T $T=29520 98400 0 0 $X=29230 $Y=98165
X214 834 1 2 58 INVD0BWP7T $T=42400 90560 0 0 $X=42110 $Y=90325
X215 846 1 2 81 INVD0BWP7T $T=47440 82720 1 0 $X=47150 $Y=78510
X216 863 1 2 805 INVD0BWP7T $T=55840 90560 1 180 $X=53870 $Y=90325
X217 867 1 2 901 INVD0BWP7T $T=79920 67040 1 0 $X=79630 $Y=62830
X218 142 1 2 903 INVD0BWP7T $T=85520 59200 0 0 $X=85230 $Y=58965
X219 151 1 2 893 INVD0BWP7T $T=85520 98400 0 0 $X=85230 $Y=98165
X220 923 1 2 912 INVD0BWP7T $T=95040 74880 0 180 $X=93070 $Y=70670
X221 239 1 2 935 INVD0BWP7T $T=110160 98400 0 180 $X=108190 $Y=94190
X222 240 1 2 951 INVD0BWP7T $T=111280 74880 0 0 $X=110990 $Y=74645
X223 948 1 2 958 INVD0BWP7T $T=111840 59200 1 0 $X=111550 $Y=54990
X224 926 1 2 969 INVD0BWP7T $T=121920 74880 0 0 $X=121630 $Y=74645
X225 978 1 2 960 INVD0BWP7T $T=126400 82720 1 180 $X=124430 $Y=82485
X226 939 1 2 955 INVD0BWP7T $T=132560 74880 0 0 $X=132270 $Y=74645
X227 217 1 2 995 INVD0BWP7T $T=139280 51360 1 180 $X=137310 $Y=51125
X228 1004 1 2 293 INVD0BWP7T $T=140960 59200 1 180 $X=138990 $Y=58965
X229 241 1 2 1011 INVD0BWP7T $T=144880 51360 0 180 $X=142910 $Y=47150
X230 184 1 2 316 INVD0BWP7T $T=146000 82720 0 0 $X=145710 $Y=82485
X231 980 1 2 1017 INVD0BWP7T $T=146560 74880 0 0 $X=146270 $Y=74645
X232 331 1 2 1012 INVD0BWP7T $T=155520 51360 0 0 $X=155230 $Y=51125
X233 229 1 2 1009 INVD0BWP7T $T=165600 106240 0 180 $X=163630 $Y=102030
X234 333 1 2 1030 INVD0BWP7T $T=166720 59200 1 180 $X=164750 $Y=58965
X235 1059 1 2 1048 INVD0BWP7T $T=176800 74880 0 180 $X=174830 $Y=70670
X236 1060 1 2 381 INVD0BWP7T $T=188560 74880 0 0 $X=188270 $Y=74645
X237 1111 1 2 1106 INVD0BWP7T $T=191920 90560 0 180 $X=189950 $Y=86350
X238 1128 1 2 399 INVD0BWP7T $T=195280 67040 0 180 $X=193310 $Y=62830
X239 411 1 2 1121 INVD0BWP7T $T=196960 82720 0 180 $X=194990 $Y=78510
X240 1071 1 2 1136 INVD0BWP7T $T=205920 82720 0 0 $X=205630 $Y=82485
X241 1081 1 2 1137 INVD0BWP7T $T=205920 98400 0 0 $X=205630 $Y=98165
X242 1160 1 2 1078 INVD0BWP7T $T=218800 59200 0 180 $X=216830 $Y=54990
X243 356 1 2 434 INVD0BWP7T $T=218240 51360 1 0 $X=217950 $Y=47150
X244 403 1 2 1166 INVD0BWP7T $T=220480 82720 0 0 $X=220190 $Y=82485
X245 1171 1 2 1113 INVD0BWP7T $T=223840 59200 1 180 $X=221870 $Y=58965
X246 419 1 2 459 INVD0BWP7T $T=228320 51360 1 0 $X=228030 $Y=47150
X247 1177 1 2 1151 INVD0BWP7T $T=230000 74880 1 180 $X=228030 $Y=74645
X248 1197 1 2 1050 INVD0BWP7T $T=241200 90560 0 180 $X=239230 $Y=86350
X249 1211 1 2 1118 INVD0BWP7T $T=256320 106240 0 180 $X=254350 $Y=102030
X250 1161 1 2 1208 INVD0BWP7T $T=259120 67040 0 0 $X=258830 $Y=66805
X251 1223 1 2 1218 INVD0BWP7T $T=270320 67040 0 180 $X=268350 $Y=62830
X252 1222 1 2 1228 INVD0BWP7T $T=275920 82720 0 0 $X=275630 $Y=82485
X253 1235 1 2 1236 INVD0BWP7T $T=292160 90560 0 0 $X=291870 $Y=90325
X254 1239 1 2 1240 INVD0BWP7T $T=295520 90560 1 0 $X=295230 $Y=86350
X255 1245 1 2 1244 INVD0BWP7T $T=307840 82720 0 180 $X=305870 $Y=78510
X256 1248 1 2 1247 INVD0BWP7T $T=309520 82720 0 180 $X=307550 $Y=78510
X257 1265 1 2 1267 INVD0BWP7T $T=339200 67040 0 0 $X=338910 $Y=66805
X258 1268 1 2 587 INVD0BWP7T $T=341440 51360 1 0 $X=341150 $Y=47150
X259 607 1 2 1256 INVD0BWP7T $T=363280 59200 0 180 $X=361310 $Y=54990
X260 614 1 2 1289 INVD0BWP7T $T=374480 82720 1 0 $X=374190 $Y=78510
X261 616 1 2 1300 INVD0BWP7T $T=380640 90560 1 0 $X=380350 $Y=86350
X262 1298 1 2 1302 INVD0BWP7T $T=381200 74880 1 0 $X=380910 $Y=70670
X263 1294 1 2 1301 INVD0BWP7T $T=383440 82720 1 0 $X=383150 $Y=78510
X264 1304 1 2 1306 INVD0BWP7T $T=386240 51360 1 180 $X=384270 $Y=51125
X265 621 1 2 1311 INVD0BWP7T $T=392960 59200 0 0 $X=392670 $Y=58965
X266 603 1 2 1314 INVD0BWP7T $T=395200 90560 0 0 $X=394910 $Y=90325
X267 1316 1 2 1312 INVD0BWP7T $T=402480 67040 0 180 $X=400510 $Y=62830
X268 664 1 2 1323 INVD0BWP7T $T=417600 74880 1 180 $X=415630 $Y=74645
X269 666 1 2 1332 INVD0BWP7T $T=419280 82720 0 0 $X=418990 $Y=82485
X270 1326 1 2 1331 INVD0BWP7T $T=420400 90560 1 0 $X=420110 $Y=86350
X271 653 1 2 1334 INVD0BWP7T $T=422080 90560 1 0 $X=421790 $Y=86350
X272 1237 513 1 2 BUFFD1P5BWP7T $T=294960 82720 1 180 $X=291870 $Y=82485
X273 1251 515 1 2 BUFFD1P5BWP7T $T=317360 59200 0 180 $X=314270 $Y=54990
X274 1258 575 1 2 BUFFD1P5BWP7T $T=336400 98400 0 180 $X=333310 $Y=94190
X275 1276 599 1 2 BUFFD1P5BWP7T $T=357680 59200 1 180 $X=354590 $Y=58965
X276 1282 635 1 2 BUFFD1P5BWP7T $T=387920 82720 1 0 $X=387630 $Y=78510
X277 725 733 1 2 BUFFD1P5BWP7T $T=461840 51360 0 0 $X=461550 $Y=51125
X278 541 1 2 546 INVD3BWP7T $T=306720 67040 0 0 $X=306430 $Y=66805
X279 560 1 2 567 INVD3BWP7T $T=319040 67040 0 0 $X=318750 $Y=66805
X280 563 1 2 569 INVD3BWP7T $T=319600 98400 1 0 $X=319310 $Y=94190
X364 860 1 2 866 BUFFD1BWP7T $T=53600 59200 1 0 $X=53310 $Y=54990
X365 866 1 2 141 BUFFD1BWP7T $T=68160 67040 1 0 $X=67870 $Y=62830
X366 915 1 2 918 BUFFD1BWP7T $T=91680 82720 0 0 $X=91390 $Y=82485
X367 924 1 2 919 BUFFD1BWP7T $T=96160 82720 1 180 $X=93630 $Y=82485
X368 986 1 2 272 BUFFD1BWP7T $T=132560 98400 0 180 $X=130030 $Y=94190
X369 1037 1 2 349 BUFFD1BWP7T $T=170640 98400 0 0 $X=170350 $Y=98165
X370 1044 1 2 345 BUFFD1BWP7T $T=173440 106240 0 180 $X=170910 $Y=102030
X371 1060 1 2 1056 BUFFD1BWP7T $T=177360 74880 1 180 $X=174830 $Y=74645
X372 1135 1 2 1110 BUFFD1BWP7T $T=208160 51360 1 180 $X=205630 $Y=51125
X373 1152 1 2 1086 BUFFD1BWP7T $T=213200 74880 0 180 $X=210670 $Y=70670
X374 482 1 2 1209 BUFFD1BWP7T $T=252400 106240 1 0 $X=252110 $Y=102030
X375 542 1 2 548 BUFFD1BWP7T $T=308400 51360 0 0 $X=308110 $Y=51125
X376 555 1 2 1250 BUFFD1BWP7T $T=313440 51360 0 0 $X=313150 $Y=51125
X377 1241 1 2 568 BUFFD1BWP7T $T=325200 82720 0 180 $X=322670 $Y=78510
X378 1301 1 2 1305 BUFFD1BWP7T $T=383440 82720 0 0 $X=383150 $Y=82485
X379 1336 1 2 681 BUFFD1BWP7T $T=432720 82720 1 180 $X=430190 $Y=82485
X380 686 1 2 1339 BUFFD1BWP7T $T=435520 106240 1 0 $X=435230 $Y=102030
X381 720 1 2 1342 BUFFD1BWP7T $T=459600 106240 1 0 $X=459310 $Y=102030
X382 734 1 2 736 BUFFD1BWP7T $T=465760 51360 0 0 $X=465470 $Y=51125
X383 1 2 DCAP4BWP7T $T=26720 82720 0 0 $X=26430 $Y=82485
X384 1 2 DCAP4BWP7T $T=48000 59200 1 0 $X=47710 $Y=54990
X385 1 2 DCAP4BWP7T $T=56960 82720 1 0 $X=56670 $Y=78510
X386 1 2 DCAP4BWP7T $T=96720 67040 0 0 $X=96430 $Y=66805
X387 1 2 DCAP4BWP7T $T=123600 51360 0 0 $X=123310 $Y=51125
X388 1 2 DCAP4BWP7T $T=141520 98400 0 0 $X=141230 $Y=98165
X389 1 2 DCAP4BWP7T $T=142080 82720 1 0 $X=141790 $Y=78510
X390 1 2 DCAP4BWP7T $T=149920 74880 1 0 $X=149630 $Y=70670
X391 1 2 DCAP4BWP7T $T=151600 82720 1 0 $X=151310 $Y=78510
X392 1 2 DCAP4BWP7T $T=161120 67040 0 0 $X=160830 $Y=66805
X393 1 2 DCAP4BWP7T $T=179040 51360 0 0 $X=178750 $Y=51125
X394 1 2 DCAP4BWP7T $T=186880 59200 0 0 $X=186590 $Y=58965
X395 1 2 DCAP4BWP7T $T=214320 98400 1 0 $X=214030 $Y=94190
X396 1 2 DCAP4BWP7T $T=221040 74880 1 0 $X=220750 $Y=70670
X397 1 2 DCAP4BWP7T $T=224400 82720 1 0 $X=224110 $Y=78510
X398 1 2 DCAP4BWP7T $T=229440 59200 0 0 $X=229150 $Y=58965
X399 1 2 DCAP4BWP7T $T=236720 74880 1 0 $X=236430 $Y=70670
X400 1 2 DCAP4BWP7T $T=237280 90560 1 0 $X=236990 $Y=86350
X401 1 2 DCAP4BWP7T $T=253520 51360 0 0 $X=253230 $Y=51125
X402 1 2 DCAP4BWP7T $T=283760 59200 0 0 $X=283470 $Y=58965
X403 1 2 DCAP4BWP7T $T=367760 74880 1 0 $X=367470 $Y=70670
X404 1 2 DCAP4BWP7T $T=371120 59200 1 0 $X=370830 $Y=54990
X405 1 2 DCAP4BWP7T $T=375600 90560 0 0 $X=375310 $Y=90325
X406 1 2 DCAP4BWP7T $T=381200 98400 0 0 $X=380910 $Y=98165
X407 1 2 DCAP4BWP7T $T=390160 98400 1 0 $X=389870 $Y=94190
X408 1 2 DCAP4BWP7T $T=399120 106240 1 0 $X=398830 $Y=102030
X409 1 2 DCAP4BWP7T $T=451760 82720 0 0 $X=451470 $Y=82485
X410 1 2 DCAP4BWP7T $T=471920 82720 0 0 $X=471630 $Y=82485
X411 1 2 DCAP4BWP7T $T=471920 106240 1 0 $X=471630 $Y=102030
X412 1 2 ICV_3 $T=35120 90560 0 0 $X=34830 $Y=90325
X413 1 2 ICV_3 $T=42400 51360 1 0 $X=42110 $Y=47150
X414 1 2 ICV_3 $T=73200 51360 0 0 $X=72910 $Y=51125
X415 1 2 ICV_3 $T=77120 74880 1 0 $X=76830 $Y=70670
X416 1 2 ICV_3 $T=87760 51360 0 0 $X=87470 $Y=51125
X417 1 2 ICV_3 $T=96160 82720 0 0 $X=95870 $Y=82485
X418 1 2 ICV_3 $T=110160 98400 0 0 $X=109870 $Y=98165
X419 1 2 ICV_3 $T=115200 90560 1 0 $X=114910 $Y=86350
X420 1 2 ICV_3 $T=119120 106240 1 0 $X=118830 $Y=102030
X421 1 2 ICV_3 $T=125840 98400 0 0 $X=125550 $Y=98165
X422 1 2 ICV_3 $T=136480 59200 0 0 $X=136190 $Y=58965
X423 1 2 ICV_3 $T=140400 51360 1 0 $X=140110 $Y=47150
X424 1 2 ICV_3 $T=146560 59200 0 0 $X=146270 $Y=58965
X425 1 2 ICV_3 $T=157200 51360 0 0 $X=156910 $Y=51125
X426 1 2 ICV_3 $T=157200 74880 0 0 $X=156910 $Y=74645
X427 1 2 ICV_3 $T=168400 51360 1 0 $X=168110 $Y=47150
X428 1 2 ICV_3 $T=171200 67040 1 0 $X=170910 $Y=62830
X429 1 2 ICV_3 $T=179040 67040 0 0 $X=178750 $Y=66805
X430 1 2 ICV_3 $T=189680 98400 0 0 $X=189390 $Y=98165
X431 1 2 ICV_3 $T=209840 106240 1 0 $X=209550 $Y=102030
X432 1 2 ICV_3 $T=214880 74880 0 0 $X=214590 $Y=74645
X433 1 2 ICV_3 $T=218800 59200 1 0 $X=218510 $Y=54990
X434 1 2 ICV_3 $T=222720 106240 1 0 $X=222430 $Y=102030
X435 1 2 ICV_3 $T=227200 51360 0 0 $X=226910 $Y=51125
X436 1 2 ICV_3 $T=241200 74880 0 0 $X=240910 $Y=74645
X437 1 2 ICV_3 $T=266960 59200 1 0 $X=266670 $Y=54990
X438 1 2 ICV_3 $T=291600 106240 1 0 $X=291310 $Y=102030
X439 1 2 ICV_3 $T=303920 82720 0 0 $X=303630 $Y=82485
X440 1 2 ICV_3 $T=308960 74880 0 0 $X=308670 $Y=74645
X441 1 2 ICV_3 $T=310640 51360 0 0 $X=310350 $Y=51125
X442 1 2 ICV_3 $T=338080 59200 0 0 $X=337790 $Y=58965
X443 1 2 ICV_3 $T=342560 98400 0 0 $X=342270 $Y=98165
X444 1 2 ICV_3 $T=357680 59200 0 0 $X=357390 $Y=58965
X445 1 2 ICV_3 $T=367200 59200 0 0 $X=366910 $Y=58965
X446 1 2 ICV_3 $T=375600 59200 0 0 $X=375310 $Y=58965
X447 1 2 ICV_3 $T=375600 106240 1 0 $X=375310 $Y=102030
X448 1 2 ICV_3 $T=385120 82720 1 0 $X=384830 $Y=78510
X449 1 2 ICV_3 $T=387360 74880 1 0 $X=387070 $Y=70670
X450 1 2 ICV_3 $T=388480 98400 0 0 $X=388190 $Y=98165
X451 1 2 ICV_3 $T=401360 74880 1 0 $X=401070 $Y=70670
X452 1 2 ICV_3 $T=409200 59200 1 0 $X=408910 $Y=54990
X453 1 2 ICV_3 $T=424320 74880 0 0 $X=424030 $Y=74645
X454 1 2 ICV_3 $T=435520 98400 0 0 $X=435230 $Y=98165
X455 1 2 ICV_3 $T=436640 59200 1 0 $X=436350 $Y=54990
X456 1 2 ICV_3 $T=438880 90560 1 0 $X=438590 $Y=86350
X457 1 2 ICV_3 $T=440560 51360 0 0 $X=440270 $Y=51125
X458 1 2 ICV_3 $T=459600 82720 0 0 $X=459310 $Y=82485
X459 1 2 ICV_3 $T=464640 82720 1 0 $X=464350 $Y=78510
X460 1 2 DCAP8BWP7T $T=23360 51360 0 0 $X=23070 $Y=51125
X461 1 2 DCAP8BWP7T $T=28960 106240 1 0 $X=28670 $Y=102030
X462 1 2 DCAP8BWP7T $T=60880 106240 1 0 $X=60590 $Y=102030
X463 1 2 DCAP8BWP7T $T=90000 67040 0 0 $X=89710 $Y=66805
X464 1 2 DCAP8BWP7T $T=98960 98400 0 0 $X=98670 $Y=98165
X465 1 2 DCAP8BWP7T $T=105680 98400 0 0 $X=105390 $Y=98165
X466 1 2 DCAP8BWP7T $T=106800 51360 1 0 $X=106510 $Y=47150
X467 1 2 DCAP8BWP7T $T=112960 51360 1 0 $X=112670 $Y=47150
X468 1 2 DCAP8BWP7T $T=119120 74880 1 0 $X=118830 $Y=70670
X469 1 2 DCAP8BWP7T $T=133680 67040 0 0 $X=133390 $Y=66805
X470 1 2 DCAP8BWP7T $T=135920 51360 1 0 $X=135630 $Y=47150
X471 1 2 DCAP8BWP7T $T=140400 90560 1 0 $X=140110 $Y=86350
X472 1 2 DCAP8BWP7T $T=152720 59200 0 0 $X=152430 $Y=58965
X473 1 2 DCAP8BWP7T $T=155520 90560 0 0 $X=155230 $Y=90325
X474 1 2 DCAP8BWP7T $T=174560 67040 0 0 $X=174270 $Y=66805
X475 1 2 DCAP8BWP7T $T=175120 90560 0 0 $X=174830 $Y=90325
X476 1 2 DCAP8BWP7T $T=177360 82720 0 0 $X=177070 $Y=82485
X477 1 2 DCAP8BWP7T $T=183520 67040 0 0 $X=183230 $Y=66805
X478 1 2 DCAP8BWP7T $T=189680 90560 0 0 $X=189390 $Y=90325
X479 1 2 DCAP8BWP7T $T=213200 67040 0 0 $X=212910 $Y=66805
X480 1 2 DCAP8BWP7T $T=214880 82720 1 0 $X=214590 $Y=78510
X481 1 2 DCAP8BWP7T $T=222720 51360 0 0 $X=222430 $Y=51125
X482 1 2 DCAP8BWP7T $T=230000 74880 0 0 $X=229710 $Y=74645
X483 1 2 DCAP8BWP7T $T=254640 98400 0 0 $X=254350 $Y=98165
X484 1 2 DCAP8BWP7T $T=258560 59200 1 0 $X=258270 $Y=54990
X485 1 2 DCAP8BWP7T $T=263600 67040 0 0 $X=263310 $Y=66805
X486 1 2 DCAP8BWP7T $T=268640 51360 0 0 $X=268350 $Y=51125
X487 1 2 DCAP8BWP7T $T=275360 74880 0 0 $X=275070 $Y=74645
X488 1 2 DCAP8BWP7T $T=278720 90560 1 0 $X=278430 $Y=86350
X489 1 2 DCAP8BWP7T $T=281520 82720 1 0 $X=281230 $Y=78510
X490 1 2 DCAP8BWP7T $T=293840 74880 0 0 $X=293550 $Y=74645
X491 1 2 DCAP8BWP7T $T=299440 59200 1 0 $X=299150 $Y=54990
X492 1 2 DCAP8BWP7T $T=299440 82720 1 0 $X=299150 $Y=78510
X493 1 2 DCAP8BWP7T $T=299440 98400 1 0 $X=299150 $Y=94190
X494 1 2 DCAP8BWP7T $T=304480 74880 0 0 $X=304190 $Y=74645
X495 1 2 DCAP8BWP7T $T=305040 74880 1 0 $X=304750 $Y=70670
X496 1 2 DCAP8BWP7T $T=313440 59200 0 0 $X=313150 $Y=58965
X497 1 2 DCAP8BWP7T $T=315680 51360 0 0 $X=315390 $Y=51125
X498 1 2 DCAP8BWP7T $T=319040 106240 1 0 $X=318750 $Y=102030
X499 1 2 DCAP8BWP7T $T=320720 67040 1 0 $X=320430 $Y=62830
X500 1 2 DCAP8BWP7T $T=321840 74880 0 0 $X=321550 $Y=74645
X501 1 2 DCAP8BWP7T $T=323520 51360 1 0 $X=323230 $Y=47150
X502 1 2 DCAP8BWP7T $T=329120 51360 0 0 $X=328830 $Y=51125
X503 1 2 DCAP8BWP7T $T=329120 98400 1 0 $X=328830 $Y=94190
X504 1 2 DCAP8BWP7T $T=338080 98400 0 0 $X=337790 $Y=98165
X505 1 2 DCAP8BWP7T $T=344800 74880 0 0 $X=344510 $Y=74645
X506 1 2 DCAP8BWP7T $T=346480 82720 1 0 $X=346190 $Y=78510
X507 1 2 DCAP8BWP7T $T=346480 98400 1 0 $X=346190 $Y=94190
X508 1 2 DCAP8BWP7T $T=353200 106240 1 0 $X=352910 $Y=102030
X509 1 2 DCAP8BWP7T $T=353760 59200 1 0 $X=353470 $Y=54990
X510 1 2 DCAP8BWP7T $T=363840 51360 1 0 $X=363550 $Y=47150
X511 1 2 DCAP8BWP7T $T=364960 51360 0 0 $X=364670 $Y=51125
X512 1 2 DCAP8BWP7T $T=365520 67040 0 0 $X=365230 $Y=66805
X513 1 2 DCAP8BWP7T $T=365520 82720 0 0 $X=365230 $Y=82485
X514 1 2 DCAP8BWP7T $T=388480 59200 0 0 $X=388190 $Y=58965
X515 1 2 DCAP8BWP7T $T=396880 74880 1 0 $X=396590 $Y=70670
X516 1 2 DCAP8BWP7T $T=404720 59200 1 0 $X=404430 $Y=54990
X517 1 2 DCAP8BWP7T $T=405840 51360 1 0 $X=405550 $Y=47150
X518 1 2 DCAP8BWP7T $T=405840 67040 0 0 $X=405550 $Y=66805
X519 1 2 DCAP8BWP7T $T=422640 90560 0 0 $X=422350 $Y=90325
X520 1 2 DCAP8BWP7T $T=424320 98400 1 0 $X=424030 $Y=94190
X521 1 2 DCAP8BWP7T $T=432160 59200 1 0 $X=431870 $Y=54990
X522 1 2 DCAP8BWP7T $T=432160 82720 1 0 $X=431870 $Y=78510
X523 1 2 DCAP8BWP7T $T=432720 82720 0 0 $X=432430 $Y=82485
X524 1 2 DCAP8BWP7T $T=433280 90560 0 0 $X=432990 $Y=90325
X525 1 2 DCAP8BWP7T $T=436080 51360 0 0 $X=435790 $Y=51125
X526 1 2 DCAP8BWP7T $T=441120 98400 0 0 $X=440830 $Y=98165
X527 1 2 DCAP8BWP7T $T=446160 67040 0 0 $X=445870 $Y=66805
X528 1 2 DCAP8BWP7T $T=446720 74880 1 0 $X=446430 $Y=70670
X529 1 2 DCAP8BWP7T $T=446720 82720 1 0 $X=446430 $Y=78510
X530 1 2 DCAP8BWP7T $T=448960 67040 1 0 $X=448670 $Y=62830
X531 1 2 DCAP8BWP7T $T=449520 74880 0 0 $X=449230 $Y=74645
X532 1 2 DCAP8BWP7T $T=455120 59200 0 0 $X=454830 $Y=58965
X533 1 2 DCAP8BWP7T $T=460160 82720 1 0 $X=459870 $Y=78510
X534 1 2 DCAP8BWP7T $T=461840 90560 1 0 $X=461550 $Y=86350
X535 1 2 DCAP8BWP7T $T=464640 82720 0 0 $X=464350 $Y=82485
X536 1 2 DCAP8BWP7T $T=466880 67040 0 0 $X=466590 $Y=66805
X537 1 2 DCAP8BWP7T $T=468000 51360 0 0 $X=467710 $Y=51125
X538 1 2 DCAP8BWP7T $T=469680 82720 1 0 $X=469390 $Y=78510
X539 2 1 DCAPBWP7T $T=21120 59200 1 0 $X=20830 $Y=54990
X540 2 1 DCAPBWP7T $T=21120 59200 0 0 $X=20830 $Y=58965
X541 2 1 DCAPBWP7T $T=21120 74880 0 0 $X=20830 $Y=74645
X542 2 1 DCAPBWP7T $T=21120 82720 0 0 $X=20830 $Y=82485
X543 2 1 DCAPBWP7T $T=21120 106240 1 0 $X=20830 $Y=102030
X544 2 1 DCAPBWP7T $T=32320 67040 0 0 $X=32030 $Y=66805
X545 2 1 DCAPBWP7T $T=41840 74880 0 0 $X=41550 $Y=74645
X546 2 1 DCAPBWP7T $T=45200 106240 1 0 $X=44910 $Y=102030
X547 2 1 DCAPBWP7T $T=45760 74880 1 0 $X=45470 $Y=70670
X548 2 1 DCAPBWP7T $T=65360 51360 1 0 $X=65070 $Y=47150
X549 2 1 DCAPBWP7T $T=65360 106240 1 0 $X=65070 $Y=102030
X550 2 1 DCAPBWP7T $T=66480 98400 1 0 $X=66190 $Y=94190
X551 2 1 DCAPBWP7T $T=74320 98400 1 0 $X=74030 $Y=94190
X552 2 1 DCAPBWP7T $T=87760 67040 1 0 $X=87470 $Y=62830
X553 2 1 DCAPBWP7T $T=91680 90560 1 0 $X=91390 $Y=86350
X554 2 1 DCAPBWP7T $T=129760 82720 0 0 $X=129470 $Y=82485
X555 2 1 DCAPBWP7T $T=129760 90560 1 0 $X=129470 $Y=86350
X556 2 1 DCAPBWP7T $T=139280 51360 0 0 $X=138990 $Y=51125
X557 2 1 DCAPBWP7T $T=144320 106240 1 0 $X=144030 $Y=102030
X558 2 1 DCAPBWP7T $T=179600 90560 0 0 $X=179310 $Y=90325
X559 2 1 DCAPBWP7T $T=182400 98400 1 0 $X=182110 $Y=94190
X560 2 1 DCAPBWP7T $T=184080 59200 1 0 $X=183790 $Y=54990
X561 2 1 DCAPBWP7T $T=185200 51360 1 0 $X=184910 $Y=47150
X562 2 1 DCAPBWP7T $T=200320 90560 0 0 $X=200030 $Y=90325
X563 2 1 DCAPBWP7T $T=211520 98400 0 0 $X=211230 $Y=98165
X564 2 1 DCAPBWP7T $T=218800 82720 0 0 $X=218510 $Y=82485
X565 2 1 DCAPBWP7T $T=221600 67040 1 0 $X=221310 $Y=62830
X566 2 1 DCAPBWP7T $T=227200 74880 1 0 $X=226910 $Y=70670
X567 2 1 DCAPBWP7T $T=258560 74880 0 0 $X=258270 $Y=74645
X568 2 1 DCAPBWP7T $T=259120 98400 1 0 $X=258830 $Y=94190
X569 2 1 DCAPBWP7T $T=265280 98400 0 0 $X=264990 $Y=98165
X570 2 1 DCAPBWP7T $T=268080 67040 0 0 $X=267790 $Y=66805
X571 2 1 DCAPBWP7T $T=272000 59200 1 0 $X=271710 $Y=54990
X572 2 1 DCAPBWP7T $T=272000 82720 1 0 $X=271710 $Y=78510
X573 2 1 DCAPBWP7T $T=273120 51360 0 0 $X=272830 $Y=51125
X574 2 1 DCAPBWP7T $T=274240 106240 1 0 $X=273950 $Y=102030
X575 2 1 DCAPBWP7T $T=277600 74880 1 0 $X=277310 $Y=70670
X576 2 1 DCAPBWP7T $T=284320 51360 0 0 $X=284030 $Y=51125
X577 2 1 DCAPBWP7T $T=291600 74880 1 0 $X=291310 $Y=70670
X578 2 1 DCAPBWP7T $T=293840 51360 1 0 $X=293550 $Y=47150
X579 2 1 DCAPBWP7T $T=306720 51360 0 0 $X=306430 $Y=51125
X580 2 1 DCAPBWP7T $T=317920 59200 0 0 $X=317630 $Y=58965
X581 2 1 DCAPBWP7T $T=326320 59200 1 0 $X=326030 $Y=54990
X582 2 1 DCAPBWP7T $T=326320 74880 0 0 $X=326030 $Y=74645
X583 2 1 DCAPBWP7T $T=326320 90560 0 0 $X=326030 $Y=90325
X584 2 1 DCAPBWP7T $T=333600 51360 0 0 $X=333310 $Y=51125
X585 2 1 DCAPBWP7T $T=349280 106240 1 0 $X=348990 $Y=102030
X586 2 1 DCAPBWP7T $T=351520 59200 0 0 $X=351230 $Y=58965
X587 2 1 DCAPBWP7T $T=352080 51360 1 0 $X=351790 $Y=47150
X588 2 1 DCAPBWP7T $T=368320 51360 1 0 $X=368030 $Y=47150
X589 2 1 DCAPBWP7T $T=377840 51360 0 0 $X=377550 $Y=51125
X590 2 1 DCAPBWP7T $T=384000 90560 0 0 $X=383710 $Y=90325
X591 2 1 DCAPBWP7T $T=389040 74880 0 0 $X=388750 $Y=74645
X592 2 1 DCAPBWP7T $T=410320 51360 1 0 $X=410030 $Y=47150
X593 2 1 DCAPBWP7T $T=410320 67040 0 0 $X=410030 $Y=66805
X594 2 1 DCAPBWP7T $T=410320 74880 1 0 $X=410030 $Y=70670
X595 2 1 DCAPBWP7T $T=417600 59200 1 0 $X=417310 $Y=54990
X596 2 1 DCAPBWP7T $T=417600 82720 0 0 $X=417310 $Y=82485
X597 2 1 DCAPBWP7T $T=422080 67040 0 0 $X=421790 $Y=66805
X598 2 1 DCAPBWP7T $T=422080 82720 1 0 $X=421790 $Y=78510
X599 2 1 DCAPBWP7T $T=428800 82720 0 0 $X=428510 $Y=82485
X600 2 1 DCAPBWP7T $T=433840 106240 1 0 $X=433550 $Y=102030
X601 2 1 DCAPBWP7T $T=437200 82720 0 0 $X=436910 $Y=82485
X602 2 1 DCAPBWP7T $T=437200 98400 1 0 $X=436910 $Y=94190
X603 2 1 DCAPBWP7T $T=452320 59200 1 0 $X=452030 $Y=54990
X604 2 1 DCAPBWP7T $T=459600 59200 1 0 $X=459310 $Y=54990
X605 2 1 DCAPBWP7T $T=461840 74880 1 0 $X=461550 $Y=70670
X606 2 1 DCAPBWP7T $T=472480 51360 1 0 $X=472190 $Y=47150
X607 2 1 DCAPBWP7T $T=472480 51360 0 0 $X=472190 $Y=51125
X608 2 1 DCAPBWP7T $T=472480 67040 1 0 $X=472190 $Y=62830
X609 1 2 ICV_4 $T=57520 51360 0 0 $X=57230 $Y=51125
X610 1 2 ICV_4 $T=72080 67040 1 0 $X=71790 $Y=62830
X611 1 2 ICV_4 $T=107360 74880 1 0 $X=107070 $Y=70670
X612 1 2 ICV_4 $T=114080 90560 0 0 $X=113790 $Y=90325
X613 1 2 ICV_4 $T=119120 51360 1 0 $X=118830 $Y=47150
X614 1 2 ICV_4 $T=156080 51360 1 0 $X=155790 $Y=47150
X615 1 2 ICV_4 $T=161120 59200 1 0 $X=160830 $Y=54990
X616 1 2 ICV_4 $T=161120 59200 0 0 $X=160830 $Y=58965
X617 1 2 ICV_4 $T=161120 67040 1 0 $X=160830 $Y=62830
X618 1 2 ICV_4 $T=161120 82720 1 0 $X=160830 $Y=78510
X619 1 2 ICV_4 $T=161120 82720 0 0 $X=160830 $Y=82485
X620 1 2 ICV_4 $T=219920 74880 0 0 $X=219630 $Y=74645
X621 1 2 ICV_4 $T=228320 106240 1 0 $X=228030 $Y=102030
X622 1 2 ICV_4 $T=230560 59200 1 0 $X=230270 $Y=54990
X623 1 2 ICV_4 $T=245120 59200 1 0 $X=244830 $Y=54990
X624 1 2 ICV_4 $T=282080 51360 1 0 $X=281790 $Y=47150
X625 1 2 ICV_4 $T=282080 82720 0 0 $X=281790 $Y=82485
X626 1 2 ICV_4 $T=282080 98400 0 0 $X=281790 $Y=98165
X627 1 2 ICV_4 $T=287120 51360 0 0 $X=286830 $Y=51125
X628 1 2 ICV_4 $T=309520 82720 1 0 $X=309230 $Y=78510
X629 1 2 ICV_4 $T=324080 90560 1 0 $X=323790 $Y=86350
X630 1 2 ICV_4 $T=351520 82720 0 0 $X=351230 $Y=82485
X631 1 2 ICV_4 $T=355440 82720 1 0 $X=355150 $Y=78510
X632 1 2 ICV_4 $T=366080 106240 1 0 $X=365790 $Y=102030
X633 1 2 ICV_4 $T=371120 51360 1 0 $X=370830 $Y=47150
X634 1 2 ICV_4 $T=408080 90560 1 0 $X=407790 $Y=86350
X635 1 2 ICV_4 $T=413120 74880 1 0 $X=412830 $Y=70670
X636 1 2 ICV_4 $T=413120 90560 1 0 $X=412830 $Y=86350
X637 1 2 ICV_4 $T=450080 51360 1 0 $X=449790 $Y=47150
X638 1 2 ICV_4 $T=450080 90560 1 0 $X=449790 $Y=86350
X639 1 2 ICV_4 $T=455120 98400 1 0 $X=454830 $Y=94190
X640 1 2 ICV_4 $T=465760 51360 1 0 $X=465470 $Y=47150
X641 537 588 539 2 1 1241 DFCNQD1BWP7T $T=346480 82720 0 180 $X=333870 $Y=78510
X642 537 647 539 2 1 1282 DFCNQD1BWP7T $T=400800 82720 1 180 $X=388190 $Y=82485
X965 1 2 ICV_8 $T=34000 51360 1 0 $X=33710 $Y=47150
X966 1 2 ICV_8 $T=76000 67040 1 0 $X=75710 $Y=62830
X967 1 2 ICV_8 $T=76000 74880 0 0 $X=75710 $Y=74645
X968 1 2 ICV_8 $T=76000 82720 0 0 $X=75710 $Y=82485
X969 1 2 ICV_8 $T=76000 106240 1 0 $X=75710 $Y=102030
X970 1 2 ICV_8 $T=118000 59200 1 0 $X=117710 $Y=54990
X971 1 2 ICV_8 $T=118000 90560 0 0 $X=117710 $Y=90325
X972 1 2 ICV_8 $T=160000 90560 1 0 $X=159710 $Y=86350
X973 1 2 ICV_8 $T=160000 90560 0 0 $X=159710 $Y=90325
X974 1 2 ICV_8 $T=202000 51360 0 0 $X=201710 $Y=51125
X975 1 2 ICV_8 $T=202000 106240 1 0 $X=201710 $Y=102030
X976 1 2 ICV_8 $T=244000 51360 1 0 $X=243710 $Y=47150
X977 1 2 ICV_8 $T=286000 51360 1 0 $X=285710 $Y=47150
X978 1 2 ICV_8 $T=286000 74880 0 0 $X=285710 $Y=74645
X979 1 2 ICV_8 $T=328000 59200 1 0 $X=327710 $Y=54990
X980 1 2 ICV_8 $T=328000 90560 1 0 $X=327710 $Y=86350
X981 1 2 ICV_8 $T=412000 82720 1 0 $X=411710 $Y=78510
X982 1 2 ICV_9 $T=20000 74880 1 0 $X=19710 $Y=70670
X983 1 2 ICV_9 $T=34000 51360 0 0 $X=33710 $Y=51125
X984 1 2 ICV_9 $T=76000 51360 0 0 $X=75710 $Y=51125
X985 1 2 ICV_9 $T=118000 90560 1 0 $X=117710 $Y=86350
X986 1 2 ICV_9 $T=160000 51360 0 0 $X=159710 $Y=51125
X987 1 2 ICV_9 $T=160000 74880 0 0 $X=159710 $Y=74645
X988 1 2 ICV_9 $T=202000 90560 1 0 $X=201710 $Y=86350
X989 1 2 ICV_9 $T=244000 74880 0 0 $X=243710 $Y=74645
X990 1 2 ICV_9 $T=286000 59200 0 0 $X=285710 $Y=58965
X991 1 2 ICV_9 $T=286000 74880 1 0 $X=285710 $Y=70670
X992 1 2 ICV_9 $T=286000 82720 1 0 $X=285710 $Y=78510
X993 1 2 ICV_9 $T=286000 82720 0 0 $X=285710 $Y=82485
X994 1 2 ICV_9 $T=286000 90560 0 0 $X=285710 $Y=90325
X995 1 2 ICV_9 $T=286000 98400 1 0 $X=285710 $Y=94190
X996 1 2 ICV_9 $T=286000 98400 0 0 $X=285710 $Y=98165
X997 1 2 ICV_9 $T=286000 106240 1 0 $X=285710 $Y=102030
X998 1 2 ICV_9 $T=328000 74880 1 0 $X=327710 $Y=70670
X999 1 2 ICV_9 $T=328000 74880 0 0 $X=327710 $Y=74645
X1000 1 2 ICV_9 $T=328000 90560 0 0 $X=327710 $Y=90325
X1001 1 2 ICV_9 $T=370000 59200 0 0 $X=369710 $Y=58965
X1002 1 2 ICV_9 $T=370000 67040 0 0 $X=369710 $Y=66805
X1003 1 2 ICV_9 $T=370000 74880 0 0 $X=369710 $Y=74645
X1004 1 2 ICV_9 $T=370000 82720 0 0 $X=369710 $Y=82485
X1005 1 2 ICV_9 $T=370000 106240 1 0 $X=369710 $Y=102030
X1006 1 2 ICV_9 $T=412000 59200 1 0 $X=411710 $Y=54990
X1007 1 2 ICV_9 $T=412000 59200 0 0 $X=411710 $Y=58965
X1008 1 2 ICV_9 $T=412000 82720 0 0 $X=411710 $Y=82485
X1009 1 2 ICV_9 $T=412000 106240 1 0 $X=411710 $Y=102030
X1010 1 2 ICV_9 $T=454000 59200 1 0 $X=453710 $Y=54990
X1011 1 2 ICV_9 $T=454000 82720 0 0 $X=453710 $Y=82485
X1012 1 2 ICV_9 $T=454000 106240 1 0 $X=453710 $Y=102030
X1054 1 2 ICV_13 $T=30640 51360 1 0 $X=30350 $Y=47150
X1055 1 2 ICV_13 $T=30640 51360 0 0 $X=30350 $Y=51125
X1056 1 2 ICV_13 $T=30640 59200 0 0 $X=30350 $Y=58965
X1057 1 2 ICV_13 $T=35120 82720 1 0 $X=34830 $Y=78510
X1058 1 2 ICV_13 $T=51920 51360 1 0 $X=51630 $Y=47150
X1059 1 2 ICV_13 $T=72640 82720 0 0 $X=72350 $Y=82485
X1060 1 2 ICV_13 $T=77120 51360 1 0 $X=76830 $Y=47150
X1061 1 2 ICV_13 $T=77120 98400 1 0 $X=76830 $Y=94190
X1062 1 2 ICV_13 $T=86640 74880 1 0 $X=86350 $Y=70670
X1063 1 2 ICV_13 $T=88320 82720 1 0 $X=88030 $Y=78510
X1064 1 2 ICV_13 $T=92240 106240 1 0 $X=91950 $Y=102030
X1065 1 2 ICV_13 $T=93360 90560 0 0 $X=93070 $Y=90325
X1066 1 2 ICV_13 $T=94480 67040 1 0 $X=94190 $Y=62830
X1067 1 2 ICV_13 $T=95040 74880 0 0 $X=94750 $Y=74645
X1068 1 2 ICV_13 $T=101760 98400 1 0 $X=101470 $Y=94190
X1069 1 2 ICV_13 $T=105120 82720 0 0 $X=104830 $Y=82485
X1070 1 2 ICV_13 $T=119120 59200 0 0 $X=118830 $Y=58965
X1071 1 2 ICV_13 $T=119120 82720 1 0 $X=118830 $Y=78510
X1072 1 2 ICV_13 $T=119120 98400 1 0 $X=118830 $Y=94190
X1073 1 2 ICV_13 $T=125280 67040 0 0 $X=124990 $Y=66805
X1074 1 2 ICV_13 $T=128080 59200 0 0 $X=127790 $Y=58965
X1075 1 2 ICV_13 $T=133120 90560 1 0 $X=132830 $Y=86350
X1076 1 2 ICV_13 $T=161120 51360 1 0 $X=160830 $Y=47150
X1077 1 2 ICV_13 $T=166160 90560 1 0 $X=165870 $Y=86350
X1078 1 2 ICV_13 $T=167840 51360 0 0 $X=167550 $Y=51125
X1079 1 2 ICV_13 $T=185760 82720 0 0 $X=185470 $Y=82485
X1080 1 2 ICV_13 $T=190240 74880 0 0 $X=189950 $Y=74645
X1081 1 2 ICV_13 $T=203120 90560 0 0 $X=202830 $Y=90325
X1082 1 2 ICV_13 $T=207600 74880 1 0 $X=207310 $Y=70670
X1083 1 2 ICV_13 $T=212640 51360 0 0 $X=212350 $Y=51125
X1084 1 2 ICV_13 $T=222160 82720 0 0 $X=221870 $Y=82485
X1085 1 2 ICV_13 $T=222720 67040 0 0 $X=222430 $Y=66805
X1086 1 2 ICV_13 $T=230000 82720 0 0 $X=229710 $Y=82485
X1087 1 2 ICV_13 $T=240640 90560 0 0 $X=240350 $Y=90325
X1088 1 2 ICV_13 $T=240640 98400 1 0 $X=240350 $Y=94190
X1089 1 2 ICV_13 $T=245120 98400 1 0 $X=244830 $Y=94190
X1090 1 2 ICV_13 $T=258560 67040 1 0 $X=258270 $Y=62830
X1091 1 2 ICV_13 $T=263040 51360 0 0 $X=262750 $Y=51125
X1092 1 2 ICV_13 $T=270880 90560 1 0 $X=270590 $Y=86350
X1093 1 2 ICV_13 $T=282640 74880 0 0 $X=282350 $Y=74645
X1094 1 2 ICV_13 $T=294960 74880 1 0 $X=294670 $Y=70670
X1095 1 2 ICV_13 $T=295520 59200 0 0 $X=295230 $Y=58965
X1096 1 2 ICV_13 $T=300560 67040 1 0 $X=300270 $Y=62830
X1097 1 2 ICV_13 $T=301120 90560 0 0 $X=300830 $Y=90325
X1098 1 2 ICV_13 $T=324640 59200 0 0 $X=324350 $Y=58965
X1099 1 2 ICV_13 $T=324640 74880 1 0 $X=324350 $Y=70670
X1100 1 2 ICV_13 $T=324640 98400 0 0 $X=324350 $Y=98165
X1101 1 2 ICV_13 $T=336400 98400 1 0 $X=336110 $Y=94190
X1102 1 2 ICV_13 $T=338080 51360 1 0 $X=337790 $Y=47150
X1103 1 2 ICV_13 $T=358240 59200 1 0 $X=357950 $Y=54990
X1104 1 2 ICV_13 $T=371120 82720 1 0 $X=370830 $Y=78510
X1105 1 2 ICV_13 $T=377280 90560 1 0 $X=376990 $Y=86350
X1106 1 2 ICV_13 $T=381200 51360 0 0 $X=380910 $Y=51125
X1107 1 2 ICV_13 $T=397440 67040 1 0 $X=397150 $Y=62830
X1108 1 2 ICV_13 $T=408640 98400 0 0 $X=408350 $Y=98165
X1109 1 2 ICV_13 $T=413120 98400 0 0 $X=412830 $Y=98165
X1110 1 2 ICV_13 $T=442800 106240 1 0 $X=442510 $Y=102030
X1111 1 2 ICV_13 $T=445600 98400 0 0 $X=445310 $Y=98165
X1112 1 2 ICV_13 $T=450640 67040 0 0 $X=450350 $Y=66805
X1113 1 2 ICV_13 $T=455120 67040 0 0 $X=454830 $Y=66805
X1114 1 2 ICV_13 $T=455120 90560 1 0 $X=454830 $Y=86350
X1115 1 2 ICV_13 $T=470800 90560 1 0 $X=470510 $Y=86350
X1116 1 2 ICV_13 $T=470800 98400 1 0 $X=470510 $Y=94190
X1117 602 604 1 1280 1287 2 IOA21D0BWP7T $T=358240 106240 1 0 $X=357950 $Y=102030
X1118 5 1 2 14 INVD1BWP7T $T=22800 59200 0 0 $X=22510 $Y=58965
X1119 13 1 2 809 INVD1BWP7T $T=26720 59200 1 180 $X=24750 $Y=58965
X1120 17 1 2 36 INVD1BWP7T $T=28960 51360 1 0 $X=28670 $Y=47150
X1121 44 1 2 82 INVD1BWP7T $T=46880 90560 1 0 $X=46590 $Y=86350
X1122 836 1 2 80 INVD1BWP7T $T=50240 59200 0 0 $X=49950 $Y=58965
X1123 31 1 2 864 INVD1BWP7T $T=51360 106240 1 0 $X=51070 $Y=102030
X1124 52 1 2 865 INVD1BWP7T $T=55840 51360 0 0 $X=55550 $Y=51125
X1125 112 1 2 53 INVD1BWP7T $T=59760 51360 0 180 $X=57790 $Y=47150
X1126 851 1 2 97 INVD1BWP7T $T=63680 59200 1 0 $X=63390 $Y=54990
X1127 830 1 2 116 INVD1BWP7T $T=64240 74880 0 0 $X=63950 $Y=74645
X1128 884 1 2 140 INVD1BWP7T $T=72080 67040 0 180 $X=70110 $Y=62830
X1129 179 1 2 175 INVD1BWP7T $T=91680 51360 0 180 $X=89710 $Y=47150
X1130 191 1 2 199 INVD1BWP7T $T=95600 82720 1 0 $X=95310 $Y=78510
X1131 928 1 2 931 INVD1BWP7T $T=96720 90560 0 0 $X=96430 $Y=90325
X1132 204 1 2 940 INVD1BWP7T $T=100080 90560 1 0 $X=99790 $Y=86350
X1133 221 1 2 933 INVD1BWP7T $T=103440 51360 0 0 $X=103150 $Y=51125
X1134 216 1 2 945 INVD1BWP7T $T=103440 59200 0 0 $X=103150 $Y=58965
X1135 949 1 2 943 INVD1BWP7T $T=110160 67040 0 0 $X=109870 $Y=66805
X1136 223 1 2 181 INVD1BWP7T $T=112960 51360 0 180 $X=110990 $Y=47150
X1137 957 1 2 950 INVD1BWP7T $T=115200 82720 0 180 $X=113230 $Y=78510
X1138 203 1 2 964 INVD1BWP7T $T=113520 82720 0 0 $X=113230 $Y=82485
X1139 232 1 2 252 INVD1BWP7T $T=124160 98400 0 0 $X=123870 $Y=98165
X1140 983 1 2 937 INVD1BWP7T $T=130320 67040 1 180 $X=128350 $Y=66805
X1141 952 1 2 936 INVD1BWP7T $T=131440 82720 0 0 $X=131150 $Y=82485
X1142 994 1 2 273 INVD1BWP7T $T=133120 90560 0 180 $X=131150 $Y=86350
X1143 993 1 2 231 INVD1BWP7T $T=138160 67040 0 0 $X=137870 $Y=66805
X1144 304 1 2 998 INVD1BWP7T $T=145440 59200 0 180 $X=143470 $Y=54990
X1145 1007 1 2 927 INVD1BWP7T $T=146000 74880 0 180 $X=144030 $Y=70670
X1146 297 1 2 975 INVD1BWP7T $T=168960 106240 1 0 $X=168670 $Y=102030
X1147 1075 1 2 1052 INVD1BWP7T $T=182400 98400 0 180 $X=180430 $Y=94190
X1148 355 1 2 1127 INVD1BWP7T $T=195280 67040 1 0 $X=194990 $Y=62830
X1149 1098 1 2 414 INVD1BWP7T $T=197520 59200 0 0 $X=197230 $Y=58965
X1150 405 1 2 1061 INVD1BWP7T $T=197520 98400 0 0 $X=197230 $Y=98165
X1151 425 1 2 418 INVD1BWP7T $T=212080 51360 1 0 $X=211790 $Y=47150
X1152 1175 1 2 452 INVD1BWP7T $T=233920 106240 0 180 $X=231950 $Y=102030
X1153 1196 1 2 1150 INVD1BWP7T $T=241200 59200 1 180 $X=239230 $Y=58965
X1154 475 1 2 1114 INVD1BWP7T $T=247920 51360 1 0 $X=247630 $Y=47150
X1155 1206 1 2 438 INVD1BWP7T $T=253520 90560 1 180 $X=251550 $Y=90325
X1156 1147 1 2 1210 INVD1BWP7T $T=256320 74880 0 180 $X=254350 $Y=70670
X1157 1200 1 2 412 INVD1BWP7T $T=257440 51360 1 180 $X=255470 $Y=51125
X1158 488 1 2 490 INVD1BWP7T $T=259120 106240 1 0 $X=258830 $Y=102030
X1159 1218 1 2 449 INVD1BWP7T $T=263600 67040 0 180 $X=261630 $Y=62830
X1160 501 1 2 1186 INVD1BWP7T $T=269200 74880 1 180 $X=267230 $Y=74645
X1161 1223 1 2 1224 INVD1BWP7T $T=272000 82720 0 180 $X=270030 $Y=78510
X1162 487 1 2 1201 INVD1BWP7T $T=275360 59200 0 180 $X=273390 $Y=54990
X1163 527 1 2 1183 INVD1BWP7T $T=292720 51360 1 180 $X=290750 $Y=51125
X1164 1233 1 2 1225 INVD1BWP7T $T=293280 74880 1 0 $X=292990 $Y=70670
X1165 1194 1 2 1227 INVD1BWP7T $T=300560 67040 0 180 $X=298590 $Y=62830
X1166 643 1 2 639 INVD1BWP7T $T=395760 98400 0 180 $X=393790 $Y=94190
X1167 1 2 ICV_14 $T=169520 59200 1 0 $X=169230 $Y=54990
X1168 1 2 ICV_14 $T=219920 98400 0 0 $X=219630 $Y=98165
X1169 1 2 ICV_14 $T=238400 51360 1 0 $X=238110 $Y=47150
X1170 1 2 ICV_14 $T=265280 82720 0 0 $X=264990 $Y=82485
X1171 1 2 ICV_14 $T=268080 74880 1 0 $X=267790 $Y=70670
X1172 1 2 ICV_14 $T=269760 98400 0 0 $X=269470 $Y=98165
X1173 1 2 ICV_14 $T=293840 98400 0 0 $X=293550 $Y=98165
X1174 1 2 ICV_14 $T=302800 59200 0 0 $X=302510 $Y=58965
X1175 1 2 ICV_14 $T=307280 106240 1 0 $X=306990 $Y=102030
X1176 1 2 ICV_14 $T=310080 67040 1 0 $X=309790 $Y=62830
X1177 1 2 ICV_14 $T=358240 98400 0 0 $X=357950 $Y=98165
X1178 1 2 ICV_14 $T=364400 74880 0 0 $X=364110 $Y=74645
X1179 1 2 ICV_14 $T=364400 82720 1 0 $X=364110 $Y=78510
X1180 1 2 ICV_14 $T=396880 90560 0 0 $X=396590 $Y=90325
X1181 1 2 ICV_14 $T=435520 74880 0 0 $X=435230 $Y=74645
X1182 1 2 ICV_14 $T=448400 106240 1 0 $X=448110 $Y=102030
X1183 1339 722 1 2 BUFFD2BWP7T $T=458480 90560 1 0 $X=458190 $Y=86350
X1184 726 732 1 2 BUFFD2BWP7T $T=462960 106240 1 0 $X=462670 $Y=102030
X1185 1342 746 1 2 BUFFD2BWP7T $T=468560 106240 1 0 $X=468270 $Y=102030
X1186 1 2 DCAP16BWP7T $T=168400 82720 0 0 $X=168110 $Y=82485
X1187 1 2 DCAP16BWP7T $T=264160 98400 1 0 $X=263870 $Y=94190
X1188 1 2 DCAP16BWP7T $T=274800 59200 0 0 $X=274510 $Y=58965
X1189 1 2 DCAP16BWP7T $T=294960 82720 0 0 $X=294670 $Y=82485
X1190 1 2 DCAP16BWP7T $T=297200 90560 1 0 $X=296910 $Y=86350
X1191 1 2 DCAP16BWP7T $T=300560 51360 1 0 $X=300270 $Y=47150
X1192 1 2 DCAP16BWP7T $T=314560 51360 1 0 $X=314270 $Y=47150
X1193 1 2 DCAP16BWP7T $T=317360 59200 1 0 $X=317070 $Y=54990
X1194 1 2 DCAP16BWP7T $T=317360 90560 0 0 $X=317070 $Y=90325
X1195 1 2 DCAP16BWP7T $T=329120 51360 1 0 $X=328830 $Y=47150
X1196 1 2 DCAP16BWP7T $T=329120 59200 0 0 $X=328830 $Y=58965
X1197 1 2 DCAP16BWP7T $T=329120 67040 0 0 $X=328830 $Y=66805
X1198 1 2 DCAP16BWP7T $T=329120 82720 0 0 $X=328830 $Y=82485
X1199 1 2 DCAP16BWP7T $T=329120 98400 0 0 $X=328830 $Y=98165
X1200 1 2 DCAP16BWP7T $T=340320 106240 1 0 $X=340030 $Y=102030
X1201 1 2 DCAP16BWP7T $T=340880 67040 0 0 $X=340590 $Y=66805
X1202 1 2 DCAP16BWP7T $T=341440 90560 0 0 $X=341150 $Y=90325
X1203 1 2 DCAP16BWP7T $T=344800 59200 1 0 $X=344510 $Y=54990
X1204 1 2 DCAP16BWP7T $T=355440 98400 1 0 $X=355150 $Y=94190
X1205 1 2 DCAP16BWP7T $T=358800 74880 1 0 $X=358510 $Y=70670
X1206 1 2 DCAP16BWP7T $T=360480 67040 1 0 $X=360190 $Y=62830
X1207 1 2 DCAP16BWP7T $T=371120 74880 1 0 $X=370830 $Y=70670
X1208 1 2 DCAP16BWP7T $T=388480 67040 1 0 $X=388190 $Y=62830
X1209 1 2 DCAP16BWP7T $T=389600 59200 1 0 $X=389310 $Y=54990
X1210 1 2 DCAP16BWP7T $T=390720 82720 1 0 $X=390430 $Y=78510
X1211 1 2 DCAP16BWP7T $T=399120 90560 1 0 $X=398830 $Y=86350
X1212 1 2 DCAP16BWP7T $T=402480 67040 1 0 $X=402190 $Y=62830
X1213 1 2 DCAP16BWP7T $T=413120 51360 0 0 $X=412830 $Y=51125
X1214 1 2 DCAP16BWP7T $T=413120 67040 1 0 $X=412830 $Y=62830
X1215 1 2 DCAP16BWP7T $T=413120 67040 0 0 $X=412830 $Y=66805
X1216 1 2 DCAP16BWP7T $T=429360 74880 1 0 $X=429070 $Y=70670
X1217 1 2 DCAP16BWP7T $T=431600 67040 1 0 $X=431310 $Y=62830
X1218 1 2 DCAP16BWP7T $T=432720 67040 0 0 $X=432430 $Y=66805
X1219 1 2 DCAP16BWP7T $T=455120 67040 1 0 $X=454830 $Y=62830
X1220 876 1 2 125 CKND1BWP7T $T=62000 74880 0 0 $X=61710 $Y=74645
X1221 171 1 2 906 CKND1BWP7T $T=88320 51360 1 0 $X=88030 $Y=47150
X1222 354 1 2 1045 CKND1BWP7T $T=175120 98400 1 180 $X=173150 $Y=98165
X1223 368 1 2 1088 CKND1BWP7T $T=185760 98400 0 180 $X=183790 $Y=94190
X1224 1178 1 2 1149 CKND1BWP7T $T=230000 82720 1 180 $X=228030 $Y=82485
X1225 433 1 2 1170 CKND1BWP7T $T=235040 51360 0 180 $X=233070 $Y=47150
X1226 512 1 2 511 CKND1BWP7T $T=275920 106240 1 0 $X=275630 $Y=102030
X1227 570 1 2 1257 CKND1BWP7T $T=322960 98400 0 0 $X=322670 $Y=98165
X1228 572 1 2 1254 CKND1BWP7T $T=323520 106240 1 0 $X=323230 $Y=102030
X1229 610 1 2 1285 CKND1BWP7T $T=365520 98400 1 0 $X=365230 $Y=94190
X1230 659 1 2 1309 CKND1BWP7T $T=417600 82720 0 180 $X=415630 $Y=78510
X1231 680 1 2 678 CKND1BWP7T $T=431040 98400 0 180 $X=429070 $Y=94190
X1232 1250 1 2 549 BUFFD3BWP7T $T=314560 51360 0 180 $X=310350 $Y=47150
X1233 661 608 1 2 BUFFD12BWP7T $T=417040 74880 1 0 $X=416750 $Y=70670
X1234 160 888 2 898 1 135 152 AOI22D1BWP7T $T=83840 106240 0 180 $X=79630 $Y=102030
X1235 1231 512 2 513 1 511 504 AOI22D1BWP7T $T=279280 98400 1 180 $X=275070 $Y=98165
X1236 524 512 2 517 1 511 519 AOI22D1BWP7T $T=281520 106240 0 180 $X=277310 $Y=102030
X1237 508 1255 2 562 1 559 566 AOI22D1BWP7T $T=321280 98400 1 180 $X=317070 $Y=98165
X1238 1261 639 2 1320 1 643 1326 AOI22D1BWP7T $T=403600 82720 0 0 $X=403310 $Y=82485
X1239 1321 639 2 1318 1 643 1325 AOI22D1BWP7T $T=404160 74880 1 0 $X=403870 $Y=70670
X1240 63 809 2 27 825 1 OAI21D1BWP7T $T=43520 74880 0 180 $X=39870 $Y=70670
X1241 633 1299 2 1303 1307 1 OAI21D1BWP7T $T=388480 98400 1 180 $X=384830 $Y=98165
X1242 661 676 1 2 BUFFD8BWP7T $T=423760 67040 0 0 $X=423470 $Y=66805
X1243 63 4 72 1 2 847 AO21D0BWP7T $T=44640 59200 0 0 $X=44350 $Y=58965
X1244 591 586 1 2 BUFFD6BWP7T $T=346480 98400 0 180 $X=339470 $Y=94190
X1245 6 4 2 1 INVD2BWP7T $T=23360 51360 1 180 $X=20830 $Y=51125
X1246 15 9 2 1 INVD2BWP7T $T=24480 98400 0 180 $X=21950 $Y=94190
X1247 76 822 2 1 INVD2BWP7T $T=48560 67040 1 180 $X=46030 $Y=66805
X1248 178 135 2 1 INVD2BWP7T $T=92240 106240 0 180 $X=89710 $Y=102030
X1249 339 917 2 1 INVD2BWP7T $T=168400 74880 1 180 $X=165870 $Y=74645
X1250 467 444 2 1 INVD2BWP7T $T=236160 82720 0 180 $X=233630 $Y=78510
X1251 1215 481 2 1 INVD2BWP7T $T=263040 82720 0 0 $X=262750 $Y=82485
X1252 1195 455 2 1 INVD2BWP7T $T=267520 90560 1 180 $X=264990 $Y=90325
X1253 1220 497 2 1 INVD2BWP7T $T=265840 51360 1 0 $X=265550 $Y=47150
X1254 499 1193 2 1 INVD2BWP7T $T=268080 74880 0 180 $X=265550 $Y=70670
X1255 1234 474 2 1 INVD2BWP7T $T=281520 74880 0 180 $X=278990 $Y=70670
X1256 1232 525 2 1 INVD2BWP7T $T=305600 59200 1 0 $X=305310 $Y=54990
X1257 568 1242 2 1 INVD2BWP7T $T=320160 74880 0 180 $X=317630 $Y=70670
X1258 708 709 2 1 INVD2BWP7T $T=446160 106240 1 0 $X=445870 $Y=102030
X1259 1335 714 2 1 INVD2BWP7T $T=448960 98400 0 0 $X=448670 $Y=98165
X1260 1337 717 2 1 INVD2BWP7T $T=457920 82720 1 0 $X=457630 $Y=78510
X1261 718 719 2 1 INVD2BWP7T $T=459040 98400 1 0 $X=458750 $Y=94190
X1262 1341 728 2 1 INVD2BWP7T $T=462400 82720 0 0 $X=462110 $Y=82485
X1263 716 730 2 1 INVD2BWP7T $T=463520 51360 1 0 $X=463230 $Y=47150
X1264 1340 739 2 1 INVD2BWP7T $T=467440 82720 1 0 $X=467150 $Y=78510
X1265 1338 741 2 1 INVD2BWP7T $T=468560 90560 1 0 $X=468270 $Y=86350
X1266 745 748 2 1 INVD2BWP7T $T=469680 82720 0 0 $X=469390 $Y=82485
X1267 550 545 1 2 1232 CKXOR2D1BWP7T $T=313440 59200 1 180 $X=308110 $Y=58965
X1268 565 571 1 2 573 CKXOR2D1BWP7T $T=320160 51360 0 0 $X=319870 $Y=51125
X1269 1279 603 1 2 1281 CKXOR2D1BWP7T $T=355440 82720 0 0 $X=355150 $Y=82485
X1270 1282 1280 1 2 601 CKXOR2D1BWP7T $T=362720 90560 1 180 $X=357390 $Y=90325
X1271 1262 1284 1 2 1279 CKXOR2D1BWP7T $T=359360 82720 1 0 $X=359070 $Y=78510
X1272 1286 1257 1 2 605 CKXOR2D1BWP7T $T=365520 82720 1 180 $X=360190 $Y=82485
X1273 617 621 1 2 1296 CKXOR2D1BWP7T $T=375600 82720 0 0 $X=375310 $Y=82485
X1274 1308 643 1 2 1317 CKXOR2D1BWP7T $T=399680 59200 1 0 $X=399390 $Y=54990
X1275 1317 653 1 2 1315 CKXOR2D1BWP7T $T=402480 90560 0 0 $X=402190 $Y=90325
X1276 516 509 505 1 2 CKXOR2D2BWP7T $T=279280 98400 0 180 $X=272830 $Y=94190
X1277 543 1243 1194 1 2 CKXOR2D2BWP7T $T=310080 67040 0 180 $X=303630 $Y=62830
X1278 680 1329 332 1 2 CKXOR2D2BWP7T $T=433280 90560 1 180 $X=426830 $Y=90325
X1279 2 1 DCAP32BWP7T $T=340880 74880 1 0 $X=340590 $Y=70670
X1280 2 1 DCAP32BWP7T $T=349280 90560 1 0 $X=348990 $Y=86350
X1281 2 1 DCAP32BWP7T $T=455120 74880 0 0 $X=454830 $Y=74645
X1282 2 1 DCAP32BWP7T $T=455120 98400 0 0 $X=454830 $Y=98165
X1283 339 343 333 228 1 2 OAI21D0BWP7T $T=168960 106240 0 180 $X=165870 $Y=102030
X1284 1110 388 1093 384 1 2 OAI21D0BWP7T $T=190800 106240 0 180 $X=187710 $Y=102030
X1285 395 1062 1118 1126 1 2 OAI21D0BWP7T $T=191360 106240 1 0 $X=191070 $Y=102030
X1286 504 1221 500 508 1 2 OAI21D0BWP7T $T=271440 106240 1 0 $X=271150 $Y=102030
X1287 519 520 522 508 1 2 OAI21D0BWP7T $T=279280 98400 0 0 $X=278990 $Y=98165
X1288 1300 1293 632 1310 1 2 OAI21D0BWP7T $T=385680 90560 0 0 $X=385390 $Y=90325
X1289 1325 1328 660 1330 1 2 OAI21D0BWP7T $T=415920 98400 1 0 $X=415630 $Y=94190
X1290 1331 1333 666 508 1 2 OAI21D0BWP7T $T=421520 98400 1 0 $X=421230 $Y=94190
X1291 515 1209 1 2 1233 XNR2D1BWP7T $T=277600 90560 0 0 $X=277310 $Y=90325
X1292 1253 512 1 2 556 XNR2D1BWP7T $T=320720 67040 0 180 $X=315390 $Y=62830
X1293 559 1256 1 2 1255 XNR2D1BWP7T $T=319600 59200 0 0 $X=319310 $Y=58965
X1294 1259 512 1 2 574 XNR2D1BWP7T $T=336960 67040 0 180 $X=331630 $Y=62830
X1295 596 1277 2 1 CKND2BWP7T $T=353200 82720 1 0 $X=352910 $Y=78510
X1296 29 1 2 810 CKND0BWP7T $T=27280 90560 0 0 $X=26990 $Y=90325
X1297 267 1 2 987 CKND0BWP7T $T=128080 98400 1 0 $X=127790 $Y=94190
X1298 274 1 2 979 CKND0BWP7T $T=152160 74880 1 0 $X=151870 $Y=70670
X1299 1079 1 2 1047 CKND0BWP7T $T=181840 67040 0 0 $X=181550 $Y=66805
X1300 1108 1 2 366 CKND0BWP7T $T=190800 59200 1 180 $X=188830 $Y=58965
X1301 409 1 2 426 CKND0BWP7T $T=226080 67040 0 0 $X=225790 $Y=66805
X1302 547 1 2 1243 CKND0BWP7T $T=309520 74880 1 0 $X=309230 $Y=70670
X1303 597 1 2 1272 CKND0BWP7T $T=353200 59200 0 0 $X=352910 $Y=58965
X1304 624 1 2 628 CKND0BWP7T $T=379520 51360 0 0 $X=379230 $Y=51125
X1305 1260 2 1257 582 1262 1264 1 AOI22D2BWP7T $T=334720 90560 0 0 $X=334430 $Y=90325
X1306 599 2 1257 595 1262 1273 1 AOI22D2BWP7T $T=357680 90560 1 180 $X=350670 $Y=90325
X1307 623 627 629 1299 1 2 MUX2ND0BWP7T $T=378400 106240 1 0 $X=378110 $Y=102030
X1308 276 1 2 991 CKBD0BWP7T $T=133120 82720 0 180 $X=130590 $Y=78510
X1309 1101 1 2 382 CKBD0BWP7T $T=189680 98400 1 180 $X=187150 $Y=98165
X1310 8 2 808 20 1 NR2D1BWP7T $T=22800 106240 1 0 $X=22510 $Y=102030
X1311 8 2 821 37 1 NR2D1BWP7T $T=28400 51360 0 0 $X=28110 $Y=51125
X1312 833 2 872 858 1 NR2D1BWP7T $T=60320 74880 0 180 $X=57790 $Y=70670
X1313 844 2 905 893 1 NR2D1BWP7T $T=83840 90560 0 0 $X=83550 $Y=90325
X1314 192 2 197 204 1 NR2D1BWP7T $T=95600 106240 1 0 $X=95310 $Y=102030
X1315 931 2 193 217 1 NR2D1BWP7T $T=100640 106240 1 0 $X=100350 $Y=102030
X1316 223 2 222 217 1 NR2D1BWP7T $T=105120 82720 1 180 $X=102590 $Y=82485
X1317 234 2 938 958 1 NR2D1BWP7T $T=110720 59200 0 0 $X=110430 $Y=58965
X1318 945 2 961 234 1 NR2D1BWP7T $T=115200 59200 1 180 $X=112670 $Y=58965
X1319 259 2 971 213 1 NR2D1BWP7T $T=121920 82720 0 0 $X=121630 $Y=82485
X1320 976 2 970 951 1 NR2D1BWP7T $T=124720 82720 0 180 $X=122190 $Y=78510
X1321 980 2 261 968 1 NR2D1BWP7T $T=126960 74880 1 180 $X=124430 $Y=74645
X1322 213 2 977 960 1 NR2D1BWP7T $T=124720 90560 0 0 $X=124430 $Y=90325
X1323 990 2 277 989 1 NR2D1BWP7T $T=134800 98400 0 180 $X=132270 $Y=94190
X1324 969 2 999 955 1 NR2D1BWP7T $T=139280 74880 1 180 $X=136750 $Y=74645
X1325 1000 2 291 294 1 NR2D1BWP7T $T=137600 67040 1 0 $X=137310 $Y=62830
X1326 317 2 294 304 1 NR2D1BWP7T $T=149360 51360 0 180 $X=146830 $Y=47150
X1327 327 2 325 1012 1 NR2D1BWP7T $T=154960 67040 0 0 $X=154670 $Y=66805
X1328 339 2 1031 332 1 NR2D1BWP7T $T=167280 82720 0 180 $X=164750 $Y=78510
X1329 1030 2 331 340 1 NR2D1BWP7T $T=167280 59200 1 0 $X=166990 $Y=54990
X1330 385 2 1059 366 1 NR2D1BWP7T $T=189120 67040 0 180 $X=186590 $Y=62830
X1331 1043 2 1075 403 1 NR2D1BWP7T $T=193040 82720 0 0 $X=192750 $Y=82485
X1332 385 2 1120 412 1 NR2D1BWP7T $T=196400 51360 0 0 $X=196110 $Y=51125
X1333 358 2 377 414 1 NR2D1BWP7T $T=214320 98400 0 180 $X=211790 $Y=94190
X1334 1113 2 1109 442 1 NR2D1BWP7T $T=219360 67040 1 0 $X=219070 $Y=62830
X1335 1169 2 1156 403 1 NR2D1BWP7T $T=223840 90560 0 180 $X=221310 $Y=86350
X1336 1174 2 448 1078 1 NR2D1BWP7T $T=225520 67040 0 180 $X=222990 $Y=62830
X1337 1216 2 1117 1208 1 NR2D1BWP7T $T=263040 106240 0 180 $X=260510 $Y=102030
X1338 1195 2 1189 1227 1 NR2D1BWP7T $T=274240 90560 1 0 $X=273950 $Y=86350
X1339 510 2 1196 1201 1 NR2D1BWP7T $T=277040 51360 1 180 $X=274510 $Y=51125
X1340 1227 2 1229 525 1 NR2D1BWP7T $T=292720 59200 0 180 $X=290190 $Y=54990
X1341 613 2 1288 598 1 NR2D1BWP7T $T=373920 98400 1 0 $X=373630 $Y=94190
X1342 376 374 1081 1061 1 2 AOI21D0BWP7T $T=184080 90560 0 180 $X=180990 $Y=86350
X1343 1159 432 1157 1061 1 2 AOI21D0BWP7T $T=215440 106240 0 180 $X=212350 $Y=102030
X1344 504 502 500 1221 1 2 AOI21D0BWP7T $T=269760 98400 1 180 $X=266670 $Y=98165
X1345 620 1291 625 626 1 2 AOI21D0BWP7T $T=378400 98400 0 0 $X=378110 $Y=98165
X1346 1300 1310 632 586 1 2 AOI21D0BWP7T $T=387360 98400 1 0 $X=387070 $Y=94190
X1347 1325 1330 660 633 1 2 AOI21D0BWP7T $T=416480 98400 0 0 $X=416190 $Y=98165
X1348 1331 1327 666 1333 1 2 AOI21D0BWP7T $T=419840 90560 0 0 $X=419550 $Y=90325
X1349 819 807 33 812 2 1 14 NR4D1BWP7T $T=31200 67040 0 180 $X=25310 $Y=62830
X1350 114 109 80 859 2 1 82 NR4D1BWP7T $T=60320 67040 1 180 $X=54430 $Y=66805
X1351 873 18 854 874 2 1 113 NR4D1BWP7T $T=55280 106240 1 0 $X=54990 $Y=102030
X1352 128 121 879 845 2 1 833 NR4D1BWP7T $T=64800 82720 1 180 $X=58910 $Y=82485
X1353 878 112 97 839 2 1 11 NR4D1BWP7T $T=65920 67040 1 180 $X=60030 $Y=66805
X1354 831 807 822 134 2 1 884 NR4D1BWP7T $T=63680 59200 0 0 $X=63390 $Y=58965
X1355 132 33 822 861 2 1 884 NR4D1BWP7T $T=65360 59200 1 0 $X=65070 $Y=54990
X1356 882 822 18 862 2 1 894 NR4D1BWP7T $T=67040 74880 0 0 $X=66750 $Y=74645
X1357 162 887 881 150 2 1 900 NR4D1BWP7T $T=85520 59200 1 180 $X=79630 $Y=58965
X1358 161 109 885 869 2 1 855 NR4D1BWP7T $T=85520 90560 0 180 $X=79630 $Y=86350
X1359 902 864 97 890 2 1 885 NR4D1BWP7T $T=82720 82720 1 0 $X=82430 $Y=78510
X1360 174 900 133 163 2 1 815 NR4D1BWP7T $T=90560 59200 0 180 $X=84670 $Y=54990
X1361 934 231 950 202 2 1 244 NR4D1BWP7T $T=105120 59200 1 0 $X=104830 $Y=54990
X1362 242 231 234 221 2 1 945 NR4D1BWP7T $T=110720 59200 1 180 $X=104830 $Y=58965
X1363 263 234 936 963 2 1 968 NR4D1BWP7T $T=128080 59200 1 180 $X=122190 $Y=58965
X1364 985 983 221 966 2 1 943 NR4D1BWP7T $T=129760 90560 0 180 $X=123870 $Y=86350
X1365 307 276 980 1023 2 1 1013 NR4D1BWP7T $T=146000 82720 1 0 $X=145710 $Y=78510
X1366 310 254 201 1025 2 1 1020 NR4D1BWP7T $T=146000 106240 1 0 $X=145710 $Y=102030
X1367 313 320 972 1015 2 1 1014 NR4D1BWP7T $T=148240 98400 1 0 $X=147950 $Y=94190
X1368 324 927 321 1031 2 1 945 NR4D1BWP7T $T=151600 74880 0 0 $X=151310 $Y=74645
X1369 326 1032 201 1021 2 1 229 NR4D1BWP7T $T=157200 106240 0 180 $X=151310 $Y=102030
X1370 362 358 356 1052 2 1 1045 NR4D1BWP7T $T=178480 98400 0 180 $X=172590 $Y=94190
X1371 1074 1078 1047 365 2 1 1064 NR4D1BWP7T $T=184080 59200 0 180 $X=178190 $Y=54990
X1372 1080 366 1056 1084 2 1 1086 NR4D1BWP7T $T=178480 74880 0 0 $X=178190 $Y=74645
X1373 1122 393 1114 1103 2 1 408 NR4D1BWP7T $T=190240 51360 1 0 $X=189950 $Y=47150
X1374 1123 1127 393 1132 2 1 399 NR4D1BWP7T $T=193040 59200 1 0 $X=192750 $Y=54990
X1375 1112 1111 403 1119 2 1 415 NR4D1BWP7T $T=193600 74880 0 0 $X=193310 $Y=74645
X1376 1092 415 1145 1130 2 1 427 NR4D1BWP7T $T=207600 67040 0 0 $X=207310 $Y=66805
X1377 424 1047 1136 1143 2 1 1141 NR4D1BWP7T $T=213200 82720 1 180 $X=207310 $Y=82485
X1378 1104 1127 1149 1153 2 1 1155 NR4D1BWP7T $T=208160 90560 1 0 $X=207870 $Y=86350
X1379 1042 428 426 1136 2 1 1111 NR4D1BWP7T $T=214880 82720 0 180 $X=208990 $Y=78510
X1380 429 425 1149 1162 2 1 1163 NR4D1BWP7T $T=213200 82720 0 0 $X=212910 $Y=82485
X1381 454 1177 456 1185 2 1 1111 NR4D1BWP7T $T=228320 82720 1 0 $X=228030 $Y=78510
X1382 1133 457 444 1185 2 1 465 NR4D1BWP7T $T=230000 98400 0 0 $X=229710 $Y=98165
X1383 1180 479 465 1198 2 1 1208 NR4D1BWP7T $T=249040 98400 0 0 $X=248750 $Y=98165
X1384 1205 436 1210 1212 2 1 442 NR4D1BWP7T $T=253520 67040 0 0 $X=253230 $Y=66805
X1385 1107 411 492 1219 2 1 1217 NR4D1BWP7T $T=259680 98400 0 0 $X=259390 $Y=98165
X1386 940 199 938 2 1 922 AN3D1BWP7T $T=102320 82720 1 180 $X=98670 $Y=82485
X1387 1061 2 347 1050 1039 1035 1 AOI31D2BWP7T $T=176240 90560 0 180 $X=169230 $Y=86350
X1388 375 2 363 1071 360 1072 1 AOI31D2BWP7T $T=181280 106240 0 180 $X=174270 $Y=102030
X1389 838 861 847 82 2 1 867 OR4D1BWP7T $T=51920 59200 0 0 $X=51630 $Y=58965
X1390 847 105 108 107 2 1 876 OR4D1BWP7T $T=56400 59200 0 0 $X=56110 $Y=58965
X1391 131 94 886 135 1 2 145 OA31D0BWP7T $T=67040 106240 1 0 $X=66750 $Y=102030
X1392 332 1030 317 949 1 2 1004 OA31D0BWP7T $T=157200 59200 0 180 $X=152430 $Y=54990
X1393 525 491 1194 518 1 2 1182 OA31D0BWP7T $T=282640 59200 0 180 $X=277870 $Y=54990
X1394 1181 2 1158 1193 481 1 AOI21D2BWP7T $T=258000 82720 0 0 $X=257710 $Y=82485
X1395 491 2 1102 1191 527 1 AOI21D2BWP7T $T=295520 51360 1 0 $X=295230 $Y=47150
X1396 3 1 5 10 2 ND2D1BWP7T $T=21680 51360 1 0 $X=21390 $Y=47150
X1397 24 1 806 21 2 ND2D1BWP7T $T=27280 98400 0 180 $X=24750 $Y=94190
X1398 27 1 804 24 2 ND2D1BWP7T $T=29520 90560 0 180 $X=26990 $Y=86350
X1399 27 1 31 19 2 ND2D1BWP7T $T=27280 98400 0 0 $X=26990 $Y=98165
X1400 3 1 35 19 2 ND2D1BWP7T $T=30640 59200 1 180 $X=28110 $Y=58965
X1401 19 1 824 55 2 ND2D1BWP7T $T=28960 74880 0 0 $X=28670 $Y=74645
X1402 27 1 43 9 2 ND2D1BWP7T $T=28960 82720 0 0 $X=28670 $Y=82485
X1403 9 1 44 41 2 ND2D1BWP7T $T=28960 90560 0 0 $X=28670 $Y=90325
X1404 4 1 47 24 2 ND2D1BWP7T $T=37920 51360 1 0 $X=37630 $Y=47150
X1405 809 1 46 21 2 ND2D1BWP7T $T=37920 59200 0 0 $X=37630 $Y=58965
X1406 50 1 812 46 2 ND2D1BWP7T $T=40160 67040 0 180 $X=37630 $Y=62830
X1407 9 1 828 21 2 ND2D1BWP7T $T=37920 74880 1 0 $X=37630 $Y=70670
X1408 9 1 829 51 2 ND2D1BWP7T $T=37920 82720 0 0 $X=37630 $Y=82485
X1409 24 1 830 55 2 ND2D1BWP7T $T=38480 82720 1 0 $X=38190 $Y=78510
X1410 24 1 834 41 2 ND2D1BWP7T $T=39040 90560 1 0 $X=38750 $Y=86350
X1411 53 1 56 832 2 ND2D1BWP7T $T=39600 98400 1 0 $X=39310 $Y=94190
X1412 21 1 50 10 2 ND2D1BWP7T $T=40160 51360 1 0 $X=39870 $Y=47150
X1413 4 1 835 36 2 ND2D1BWP7T $T=40160 51360 0 0 $X=39870 $Y=51125
X1414 63 1 836 55 2 ND2D1BWP7T $T=42960 67040 0 180 $X=40430 $Y=62830
X1415 9 1 62 55 2 ND2D1BWP7T $T=41280 59200 1 0 $X=40990 $Y=54990
X1416 63 1 61 59 2 ND2D1BWP7T $T=44080 98400 0 180 $X=41550 $Y=94190
X1417 824 1 839 66 2 ND2D1BWP7T $T=42960 67040 1 0 $X=42670 $Y=62830
X1418 809 1 840 69 2 ND2D1BWP7T $T=42960 82720 1 0 $X=42670 $Y=78510
X1419 55 1 67 10 2 ND2D1BWP7T $T=45760 59200 0 180 $X=43230 $Y=54990
X1420 63 1 827 3 2 ND2D1BWP7T $T=44640 51360 0 0 $X=44350 $Y=51125
X1421 36 1 73 55 2 ND2D1BWP7T $T=47440 51360 0 180 $X=44910 $Y=47150
X1422 4 1 846 19 2 ND2D1BWP7T $T=45760 59200 1 0 $X=45470 $Y=54990
X1423 3 1 851 36 2 ND2D1BWP7T $T=47440 51360 1 0 $X=47150 $Y=47150
X1424 19 1 79 21 2 ND2D1BWP7T $T=48000 59200 0 0 $X=47710 $Y=58965
X1425 90 1 837 83 2 ND2D1BWP7T $T=51920 51360 0 180 $X=49390 $Y=47150
X1426 96 1 859 865 2 ND2D1BWP7T $T=53600 51360 0 0 $X=53310 $Y=51125
X1427 35 1 103 828 2 ND2D1BWP7T $T=54160 74880 1 0 $X=53870 $Y=70670
X1428 851 1 861 60 2 ND2D1BWP7T $T=63680 59200 0 180 $X=61150 $Y=54990
X1429 124 1 879 849 2 ND2D1BWP7T $T=63680 74880 0 180 $X=61150 $Y=70670
X1430 124 1 110 79 2 ND2D1BWP7T $T=69280 51360 0 180 $X=66750 $Y=47150
X1431 846 1 884 142 2 ND2D1BWP7T $T=73200 59200 0 180 $X=70670 $Y=54990
X1432 124 1 892 828 2 ND2D1BWP7T $T=70960 74880 1 0 $X=70670 $Y=70670
X1433 840 1 894 143 2 ND2D1BWP7T $T=82160 74880 1 180 $X=79630 $Y=74645
X1434 143 1 121 902 2 ND2D1BWP7T $T=79920 82720 1 0 $X=79630 $Y=78510
X1435 180 1 911 910 2 ND2D1BWP7T $T=92240 59200 1 180 $X=89710 $Y=58965
X1436 177 1 913 182 2 ND2D1BWP7T $T=90560 51360 0 0 $X=90270 $Y=51125
X1437 177 1 183 180 2 ND2D1BWP7T $T=93920 59200 0 180 $X=91390 $Y=54990
X1438 177 1 188 200 2 ND2D1BWP7T $T=92800 51360 0 0 $X=92510 $Y=51125
X1439 910 1 920 185 2 ND2D1BWP7T $T=92800 59200 0 0 $X=92510 $Y=58965
X1440 177 1 926 917 2 ND2D1BWP7T $T=94480 67040 0 0 $X=94190 $Y=66805
X1441 187 1 195 198 2 ND2D1BWP7T $T=95040 59200 1 0 $X=94750 $Y=54990
X1442 200 1 194 910 2 ND2D1BWP7T $T=97840 51360 0 180 $X=95310 $Y=47150
X1443 200 1 207 198 2 ND2D1BWP7T $T=97280 59200 1 0 $X=96990 $Y=54990
X1444 182 1 923 198 2 ND2D1BWP7T $T=101760 51360 0 180 $X=99230 $Y=47150
X1445 214 1 209 910 2 ND2D1BWP7T $T=101760 59200 0 180 $X=99230 $Y=54990
X1446 198 1 939 185 2 ND2D1BWP7T $T=100640 51360 0 0 $X=100350 $Y=51125
X1447 220 1 928 200 2 ND2D1BWP7T $T=104000 51360 0 180 $X=101470 $Y=47150
X1448 214 1 216 198 2 ND2D1BWP7T $T=104000 59200 0 180 $X=101470 $Y=54990
X1449 199 1 942 940 2 ND2D1BWP7T $T=102320 90560 1 0 $X=102030 $Y=86350
X1450 911 1 946 935 2 ND2D1BWP7T $T=103440 98400 0 0 $X=103150 $Y=98165
X1451 182 1 948 220 2 ND2D1BWP7T $T=104560 51360 1 0 $X=104270 $Y=47150
X1452 948 1 230 179 2 ND2D1BWP7T $T=105120 51360 0 0 $X=104830 $Y=51125
X1453 209 1 947 937 2 ND2D1BWP7T $T=107360 74880 0 180 $X=104830 $Y=70670
X1454 179 1 235 237 2 ND2D1BWP7T $T=107920 67040 0 0 $X=107630 $Y=66805
X1455 218 1 254 967 2 ND2D1BWP7T $T=112960 98400 0 0 $X=112670 $Y=98165
X1456 187 1 247 264 2 ND2D1BWP7T $T=121920 59200 1 0 $X=121630 $Y=54990
X1457 923 1 968 269 2 ND2D1BWP7T $T=125840 51360 0 0 $X=125550 $Y=51125
X1458 270 1 981 264 2 ND2D1BWP7T $T=129760 59200 0 180 $X=127230 $Y=54990
X1459 212 1 980 957 2 ND2D1BWP7T $T=128640 82720 1 0 $X=128350 $Y=78510
X1460 993 1 989 237 2 ND2D1BWP7T $T=132560 74880 0 180 $X=130030 $Y=70670
X1461 187 1 949 910 2 ND2D1BWP7T $T=131440 59200 0 0 $X=131150 $Y=58965
X1462 985 1 280 279 2 ND2D1BWP7T $T=132560 90560 0 0 $X=132270 $Y=90325
X1463 187 1 978 998 2 ND2D1BWP7T $T=134240 59200 0 0 $X=133950 $Y=58965
X1464 998 1 957 180 2 ND2D1BWP7T $T=139840 59200 0 180 $X=137310 $Y=54990
X1465 264 1 292 214 2 ND2D1BWP7T $T=139840 59200 1 0 $X=139550 $Y=54990
X1466 295 1 993 917 2 ND2D1BWP7T $T=139840 67040 0 0 $X=139550 $Y=66805
X1467 994 1 966 1007 2 ND2D1BWP7T $T=139840 90560 0 0 $X=139550 $Y=90325
X1468 180 1 232 264 2 ND2D1BWP7T $T=140960 51360 0 0 $X=140670 $Y=51125
X1469 998 1 994 270 2 ND2D1BWP7T $T=144320 67040 0 180 $X=141790 $Y=62830
X1470 270 1 984 910 2 ND2D1BWP7T $T=144320 59200 0 0 $X=144030 $Y=58965
X1471 998 1 1008 214 2 ND2D1BWP7T $T=146560 67040 0 180 $X=144030 $Y=62830
X1472 182 1 1007 910 2 ND2D1BWP7T $T=145440 67040 0 0 $X=145150 $Y=66805
X1473 220 1 251 185 2 ND2D1BWP7T $T=157200 74880 0 180 $X=154670 $Y=70670
X1474 910 1 1028 917 2 ND2D1BWP7T $T=163920 90560 1 0 $X=163630 $Y=86350
X1475 251 1 1020 1028 2 ND2D1BWP7T $T=166160 98400 0 180 $X=163630 $Y=94190
X1476 333 1 1024 340 2 ND2D1BWP7T $T=165040 59200 1 0 $X=164750 $Y=54990
X1477 341 1 317 322 2 ND2D1BWP7T $T=167840 51360 1 180 $X=165310 $Y=51125
X1478 998 1 338 185 2 ND2D1BWP7T $T=169520 82720 0 180 $X=166990 $Y=78510
X1479 1058 1 1077 1079 2 ND2D1BWP7T $T=180720 67040 1 0 $X=180430 $Y=62830
X1480 1058 1 1116 404 2 ND2D1BWP7T $T=197520 59200 1 180 $X=194990 $Y=58965
X1481 1108 1 1163 1165 2 ND2D1BWP7T $T=217680 74880 0 0 $X=217390 $Y=74645
X1482 1173 1 1172 1040 2 ND2D1BWP7T $T=226640 90560 0 180 $X=224110 $Y=86350
X1483 435 1 1169 1175 2 ND2D1BWP7T $T=225520 82720 0 0 $X=225230 $Y=82485
X1484 1140 1 1065 445 2 ND2D1BWP7T $T=228320 51360 0 180 $X=225790 $Y=47150
X1485 449 1 379 455 2 ND2D1BWP7T $T=226080 59200 1 0 $X=225790 $Y=54990
X1486 458 1 1108 455 2 ND2D1BWP7T $T=230560 59200 0 180 $X=228030 $Y=54990
X1487 458 1 355 461 2 ND2D1BWP7T $T=230000 51360 0 0 $X=229710 $Y=51125
X1488 1183 1 423 1186 2 ND2D1BWP7T $T=231680 59200 0 0 $X=231390 $Y=58965
X1489 1183 1 462 461 2 ND2D1BWP7T $T=235040 51360 1 180 $X=232510 $Y=51125
X1490 1186 1 1098 449 2 ND2D1BWP7T $T=235040 67040 0 180 $X=232510 $Y=62830
X1491 463 1 1164 1179 2 ND2D1BWP7T $T=235040 90560 0 180 $X=232510 $Y=86350
X1492 1183 1 1160 455 2 ND2D1BWP7T $T=236720 59200 0 180 $X=234190 $Y=54990
X1493 463 1 468 1073 2 ND2D1BWP7T $T=237280 90560 0 180 $X=234750 $Y=86350
X1494 472 1 1058 455 2 ND2D1BWP7T $T=238400 59200 1 180 $X=235870 $Y=58965
X1495 472 1 467 1193 2 ND2D1BWP7T $T=238400 59200 1 0 $X=238110 $Y=54990
X1496 474 1 1040 1186 2 ND2D1BWP7T $T=241200 74880 0 180 $X=238670 $Y=70670
X1497 1200 1 372 1204 2 ND2D1BWP7T $T=249040 59200 1 0 $X=248750 $Y=54990
X1498 478 1 1175 483 2 ND2D1BWP7T $T=249600 82720 0 0 $X=249310 $Y=82485
X1499 481 1 1206 478 2 ND2D1BWP7T $T=250720 74880 0 0 $X=250430 $Y=74645
X1500 483 1 1188 1193 2 ND2D1BWP7T $T=254080 82720 1 180 $X=251550 $Y=82485
X1501 483 1 419 455 2 ND2D1BWP7T $T=255760 90560 1 180 $X=253230 $Y=90325
X1502 481 1 1200 487 2 ND2D1BWP7T $T=258560 59200 0 180 $X=256030 $Y=54990
X1503 474 1 1173 455 2 ND2D1BWP7T $T=256320 90560 0 0 $X=256030 $Y=90325
X1504 474 1 1147 1193 2 ND2D1BWP7T $T=259120 74880 0 180 $X=256590 $Y=70670
X1505 489 1 1198 484 2 ND2D1BWP7T $T=260240 59200 1 180 $X=257710 $Y=58965
X1506 472 1 1171 487 2 ND2D1BWP7T $T=260800 51360 1 180 $X=258270 $Y=51125
X1507 475 1 1217 489 2 ND2D1BWP7T $T=260240 51360 1 0 $X=259950 $Y=47150
X1508 1183 1 475 487 2 ND2D1BWP7T $T=263040 51360 1 180 $X=260510 $Y=51125
X1509 494 1 1161 483 2 ND2D1BWP7T $T=263600 67040 1 180 $X=261070 $Y=66805
X1510 472 1 1140 461 2 ND2D1BWP7T $T=265840 51360 0 180 $X=263310 $Y=47150
X1511 1193 1 447 458 2 ND2D1BWP7T $T=266960 59200 0 180 $X=264430 $Y=54990
X1512 1183 1 1220 1193 2 ND2D1BWP7T $T=268640 51360 1 180 $X=266110 $Y=51125
X1513 487 1 498 458 2 ND2D1BWP7T $T=272000 59200 0 180 $X=269470 $Y=54990
X1514 431 1 408 1226 2 ND2D1BWP7T $T=272560 51360 1 0 $X=272270 $Y=47150
X1515 494 1 1096 496 2 ND2D1BWP7T $T=274800 59200 1 180 $X=272270 $Y=58965
X1516 1229 1 1203 487 2 ND2D1BWP7T $T=278160 59200 0 180 $X=275630 $Y=54990
X1517 493 1 507 514 2 ND2D1BWP7T $T=279840 51360 1 180 $X=277310 $Y=51125
X1518 494 1 1079 474 2 ND2D1BWP7T $T=280960 67040 1 0 $X=280670 $Y=62830
X1519 1233 1 1192 1227 2 ND2D1BWP7T $T=292720 67040 1 180 $X=290190 $Y=66805
X1520 525 1 1191 1225 2 ND2D1BWP7T $T=298880 67040 0 180 $X=296350 $Y=62830
X1521 5 1 804 17 2 803 22 OAI211D1BWP7T $T=22800 74880 0 0 $X=22510 $Y=74645
X1522 35 1 30 15 2 32 22 OAI211D1BWP7T $T=28960 106240 0 180 $X=25310 $Y=102030
X1523 42 1 819 7 2 34 28 OAI211D1BWP7T $T=30640 82720 0 180 $X=26990 $Y=78510
X1524 827 1 84 6 2 857 8 OAI211D1BWP7T $T=48560 51360 0 0 $X=48270 $Y=51125
X1525 117 1 865 111 2 874 20 OAI211D1BWP7T $T=61440 98400 1 180 $X=57790 $Y=98165
X1526 827 1 84 6 2 120 8 OAI211D1BWP7T $T=61440 51360 0 0 $X=61150 $Y=51125
X1527 827 1 84 6 2 887 8 OAI211D1BWP7T $T=68720 51360 1 180 $X=65070 $Y=51125
X1528 299 1 999 1012 2 1013 308 OAI211D1BWP7T $T=143200 74880 0 0 $X=142910 $Y=74645
X1529 984 1 1017 319 2 1027 1024 OAI211D1BWP7T $T=149360 59200 0 0 $X=149070 $Y=58965
X1530 1033 1 941 1024 2 982 327 OAI211D1BWP7T $T=157200 67040 0 180 $X=153550 $Y=62830
X1531 1008 1 979 314 2 1032 336 OAI211D1BWP7T $T=168400 67040 1 180 $X=164750 $Y=66805
X1532 419 1 1128 1191 2 471 1195 OAI211D1BWP7T $T=237280 90560 0 0 $X=236990 $Y=90325
X1533 1173 1 1187 1192 2 1168 1195 OAI211D1BWP7T $T=237280 98400 1 0 $X=236990 $Y=94190
X1534 1200 1 1073 1201 2 1143 1192 OAI211D1BWP7T $T=251840 82720 0 180 $X=248190 $Y=78510
X1535 1171 1 1139 491 2 1216 1192 OAI211D1BWP7T $T=260240 59200 0 0 $X=259950 $Y=58965
X1536 1173 1 1206 1215 2 1219 499 OAI211D1BWP7T $T=260800 98400 1 0 $X=260510 $Y=94190
X1537 498 1 1140 503 2 1212 1215 OAI211D1BWP7T $T=267520 59200 0 0 $X=267230 $Y=58965
X1538 1293 1 1290 616 2 1258 609 OAI211D1BWP7T $T=377280 90560 0 180 $X=373630 $Y=86350
X1539 116 2 88 892 891 1 820 NR4D2BWP7T $T=95040 74880 1 180 $X=81870 $Y=74645
X1540 956 2 944 274 936 1 265 NR4D2BWP7T $T=123040 51360 1 0 $X=122750 $Y=47150
X1541 438 2 412 473 1 NR2XD0BWP7T $T=254640 51360 1 0 $X=254350 $Y=47150
X1542 1210 2 1038 485 1 NR2XD0BWP7T $T=255760 59200 0 0 $X=255470 $Y=58965
X1543 1208 2 495 477 1 NR2XD0BWP7T $T=262480 74880 1 0 $X=262190 $Y=70670
X1544 823 1 811 831 54 48 2 ND4D1BWP7T $T=37920 98400 0 0 $X=37630 $Y=98165
X1545 829 1 43 804 65 841 2 ND4D1BWP7T $T=41280 90560 1 0 $X=40990 $Y=86350
X1546 836 1 64 66 71 844 2 ND4D1BWP7T $T=42400 67040 0 0 $X=42110 $Y=66805
X1547 840 1 53 47 850 74 2 ND4D1BWP7T $T=45200 98400 0 0 $X=44910 $Y=98165
X1548 76 1 43 828 64 854 2 ND4D1BWP7T $T=46880 82720 0 0 $X=46590 $Y=82485
X1549 840 1 87 92 79 89 2 ND4D1BWP7T $T=50240 74880 0 0 $X=49950 $Y=74645
X1550 16 1 865 863 818 871 2 ND4D1BWP7T $T=60320 90560 0 180 $X=56110 $Y=86350
X1551 846 1 148 811 827 890 2 ND4D1BWP7T $T=73200 51360 0 180 $X=68990 $Y=47150
X1552 836 1 142 144 147 146 2 ND4D1BWP7T $T=69280 59200 0 0 $X=68990 $Y=58965
X1553 117 1 811 848 825 149 2 ND4D1BWP7T $T=69280 67040 0 0 $X=68990 $Y=66805
X1554 840 1 143 73 144 900 2 ND4D1BWP7T $T=79920 59200 1 0 $X=79630 $Y=54990
X1555 181 1 913 919 922 189 2 ND4D1BWP7T $T=91680 82720 1 0 $X=91390 $Y=78510
X1556 926 1 933 935 932 215 2 ND4D1BWP7T $T=97840 98400 1 0 $X=97550 $Y=94190
X1557 194 1 184 933 240 956 2 ND4D1BWP7T $T=107360 51360 0 0 $X=107070 $Y=51125
X1558 948 1 957 954 222 238 2 ND4D1BWP7T $T=113520 82720 0 180 $X=109310 $Y=78510
X1559 246 1 937 248 237 256 2 ND4D1BWP7T $T=111280 74880 1 0 $X=110990 $Y=70670
X1560 267 1 975 938 921 260 2 ND4D1BWP7T $T=126400 98400 0 180 $X=122190 $Y=94190
X1561 939 1 248 978 993 285 2 ND4D1BWP7T $T=132560 74880 1 0 $X=132270 $Y=70670
X1562 994 1 979 226 288 286 2 ND4D1BWP7T $T=140400 90560 0 180 $X=136190 $Y=86350
X1563 984 1 979 237 1005 296 2 ND4D1BWP7T $T=143200 74880 1 180 $X=138990 $Y=74645
X1564 226 1 1008 184 1007 302 2 ND4D1BWP7T $T=142080 82720 0 0 $X=141790 $Y=82485
X1565 952 1 292 965 241 1014 2 ND4D1BWP7T $T=142080 90560 0 0 $X=141790 $Y=90325
X1566 1151 1 1150 1147 420 1095 2 ND4D1BWP7T $T=212640 59200 0 180 $X=208430 $Y=54990
X1567 435 1 355 418 1158 1103 2 ND4D1BWP7T $T=218240 67040 0 180 $X=214030 $Y=62830
X1568 1040 1 1108 430 434 1146 2 ND4D1BWP7T $T=221040 59200 1 180 $X=216830 $Y=58965
X1569 1171 1 447 379 1151 1041 2 ND4D1BWP7T $T=225520 59200 0 180 $X=221310 $Y=54990
X1570 1161 1 443 1150 1170 1134 2 ND4D1BWP7T $T=227200 74880 0 180 $X=222990 $Y=70670
X1571 1166 1 355 460 1179 1060 2 ND4D1BWP7T $T=228880 67040 1 0 $X=228590 $Y=62830
X1572 462 1 1175 1182 448 1084 2 ND4D1BWP7T $T=232800 74880 0 180 $X=228590 $Y=70670
X1573 467 1 462 1188 1170 1167 2 ND4D1BWP7T $T=236720 74880 0 180 $X=232510 $Y=70670
X1574 1203 1 409 1147 477 476 2 ND4D1BWP7T $T=251840 74880 0 180 $X=247630 $Y=70670
X1575 1206 1 404 1202 1117 1099 2 ND4D1BWP7T $T=252400 98400 0 180 $X=248190 $Y=94190
X1576 841 121 157 904 160 1 2 OAI31D1BWP7T $T=81600 98400 0 0 $X=81310 $Y=98165
X1577 1045 1076 373 1085 368 1 2 OAI31D1BWP7T $T=180720 98400 0 0 $X=180430 $Y=98165
X1578 1141 417 1100 1129 405 1 2 OAI31D1BWP7T $T=209840 106240 0 180 $X=205630 $Y=102030
X1579 1137 1138 1097 1144 368 1 2 OAI31D1BWP7T $T=207600 98400 0 0 $X=207310 $Y=98165
X1580 1232 1227 1230 1195 1228 1 2 OAI31D1BWP7T $T=282080 82720 1 180 $X=277870 $Y=82485
X1581 873 906 901 164 169 1 2 AOI31D0BWP7T $T=84400 106240 1 0 $X=84110 $Y=102030
X1582 1123 1105 1117 396 1088 1 2 AOI31D0BWP7T $T=194720 98400 0 180 $X=191070 $Y=94190
X1583 413 410 1131 407 395 1 2 AOI31D0BWP7T $T=198640 106240 0 180 $X=194990 $Y=102030
X1584 835 1 16 819 2 838 ND3D0BWP7T $T=41840 59200 0 0 $X=41550 $Y=58965
X1585 75 1 76 44 2 855 ND3D0BWP7T $T=46880 106240 1 0 $X=46590 $Y=102030
X1586 64 1 87 853 2 858 ND3D0BWP7T $T=48560 67040 0 0 $X=48270 $Y=66805
X1587 67 1 806 65 2 94 ND3D0BWP7T $T=50240 90560 1 0 $X=49950 $Y=86350
X1588 865 1 62 73 2 104 ND3D0BWP7T $T=55280 51360 1 0 $X=54990 $Y=47150
X1589 60 1 16 865 2 122 ND3D0BWP7T $T=60320 98400 1 0 $X=60030 $Y=94190
X1590 877 1 872 132 2 886 ND3D0BWP7T $T=65920 67040 0 0 $X=65630 $Y=66805
X1591 897 1 896 147 2 155 ND3D0BWP7T $T=79920 74880 1 0 $X=79630 $Y=70670
X1592 939 1 934 922 2 914 ND3D0BWP7T $T=101200 74880 1 180 $X=98110 $Y=74645
X1593 992 1 973 941 2 278 ND3D0BWP7T $T=131440 67040 1 0 $X=131150 $Y=62830
X1594 1016 1 964 309 2 1015 ND3D0BWP7T $T=148240 98400 0 180 $X=145150 $Y=94190
X1595 232 1 1034 1029 2 328 ND3D0BWP7T $T=156640 90560 0 180 $X=153550 $Y=86350
X1596 1058 1 351 355 2 1051 ND3D0BWP7T $T=176800 67040 0 180 $X=173710 $Y=62830
X1597 379 1 1098 380 2 1082 ND3D0BWP7T $T=188560 59200 0 180 $X=185470 $Y=54990
X1598 1112 1 1066 1109 2 1046 ND3D0BWP7T $T=192480 67040 1 180 $X=189390 $Y=66805
X1599 1161 1 1147 431 2 401 ND3D0BWP7T $T=221040 74880 0 180 $X=217950 $Y=70670
X1600 1220 1 431 1140 2 1214 ND3D0BWP7T $T=267520 67040 0 180 $X=264430 $Y=62830
X1601 816 1 2 842 81 856 86 NR4D0BWP7T $T=53040 98400 1 180 $X=49390 $Y=98165
X1602 821 1 2 14 80 860 95 NR4D0BWP7T $T=50240 59200 1 0 $X=49950 $Y=54990
X1603 805 1 2 80 86 875 115 NR4D0BWP7T $T=56960 98400 1 0 $X=56670 $Y=94190
X1604 881 1 2 11 108 877 72 NR4D0BWP7T $T=62560 67040 0 180 $X=58910 $Y=62830
X1605 889 1 2 26 25 895 893 NR4D0BWP7T $T=69840 90560 0 0 $X=69550 $Y=90325
X1606 88 1 2 881 26 896 903 NR4D0BWP7T $T=79920 67040 0 0 $X=79630 $Y=66805
X1607 158 1 2 103 116 897 864 NR4D0BWP7T $T=83280 74880 1 0 $X=82990 $Y=70670
X1608 916 1 2 914 912 915 175 NR4D0BWP7T $T=93360 74880 0 180 $X=89710 $Y=70670
X1609 202 1 2 191 927 929 912 NR4D0BWP7T $T=98400 74880 0 180 $X=94750 $Y=70670
X1610 233 1 2 944 186 924 225 NR4D0BWP7T $T=107920 90560 0 180 $X=104270 $Y=86350
X1611 947 1 2 943 951 954 955 NR4D0BWP7T $T=106800 74880 0 0 $X=106510 $Y=74645
X1612 959 1 2 225 223 953 221 NR4D0BWP7T $T=111840 82720 1 180 $X=108190 $Y=82485
X1613 966 1 2 253 250 255 950 NR4D0BWP7T $T=115200 106240 0 180 $X=111550 $Y=102030
X1614 943 1 2 258 239 973 927 NR4D0BWP7T $T=125280 67040 1 180 $X=121630 $Y=66805
X1615 966 1 2 252 931 974 258 NR4D0BWP7T $T=125280 106240 0 180 $X=121630 $Y=102030
X1616 211 1 2 989 987 271 252 NR4D0BWP7T $T=128640 98400 0 0 $X=128350 $Y=98165
X1617 274 1 2 275 958 992 231 NR4D0BWP7T $T=133120 59200 0 180 $X=129470 $Y=54990
X1618 281 1 2 946 987 996 273 NR4D0BWP7T $T=134240 106240 0 180 $X=130590 $Y=102030
X1619 230 1 2 968 283 1001 275 NR4D0BWP7T $T=133680 59200 1 0 $X=133390 $Y=54990
X1620 297 1 2 946 204 1006 289 NR4D0BWP7T $T=141520 98400 1 180 $X=137870 $Y=98165
X1621 321 1 2 274 320 1018 325 NR4D0BWP7T $T=150480 90560 1 0 $X=150190 $Y=86350
X1622 1026 1 2 1020 1014 323 201 NR4D0BWP7T $T=151600 98400 0 0 $X=151310 $Y=98165
X1623 1046 1 2 1057 359 1063 1065 NR4D0BWP7T $T=175120 59200 1 0 $X=174830 $Y=54990
X1624 1119 1 2 1113 1043 1089 390 NR4D0BWP7T $T=193600 74880 0 180 $X=189950 $Y=70670
X1625 1172 1 2 1169 1052 1157 438 NR4D0BWP7T $T=226080 98400 0 180 $X=222430 $Y=94190
X1626 426 1 2 444 358 1187 390 NR4D0BWP7T $T=231120 98400 1 0 $X=230830 $Y=94190
X1627 466 1 2 468 436 469 1189 NR4D0BWP7T $T=235040 106240 1 0 $X=234750 $Y=102030
X1628 1134 1043 2 1071 1 NR2D2BWP7T $T=199200 82720 1 180 $X=194990 $Y=82485
X1629 240 247 926 226 2 1 965 AN4D1BWP7T $T=111280 90560 1 0 $X=110990 $Y=86350
X1630 964 299 1006 301 2 1 305 AN4D1BWP7T $T=141520 98400 1 0 $X=141230 $Y=94190
X1631 1140 431 430 1150 2 1 1069 AN4D1BWP7T $T=215440 59200 1 180 $X=211230 $Y=58965
X1632 473 1190 1160 470 2 1 1178 AN4D1BWP7T $T=240080 51360 1 180 $X=235870 $Y=51125
X1633 1207 485 1200 484 2 1 354 AN4D1BWP7T $T=255760 59200 1 180 $X=251550 $Y=58965
X1634 1205 1 2 1184 BUFFD0BWP7T $T=251280 67040 0 0 $X=250990 $Y=66805
X1635 519 1 2 528 BUFFD0BWP7T $T=291600 98400 0 0 $X=291310 $Y=98165
X1636 895 166 168 907 169 2 1 AOI31D1BWP7T $T=85520 90560 1 0 $X=85230 $Y=86350
X1637 170 909 172 176 178 2 1 AOI31D1BWP7T $T=87760 98400 0 0 $X=87470 $Y=98165
X1638 334 910 1029 329 302 2 1 AOI31D1BWP7T $T=157200 82720 1 180 $X=152990 $Y=82485
X1639 1079 1083 369 1089 1088 2 1 AOI31D1BWP7T $T=181840 74880 1 0 $X=181550 $Y=70670
X1640 1096 379 1068 1063 375 2 1 AOI31D1BWP7T $T=186880 67040 0 180 $X=182670 $Y=62830
X1641 1074 1105 387 1107 1088 2 1 AOI31D1BWP7T $T=187440 98400 1 0 $X=187150 $Y=94190
X1642 397 394 392 1066 375 2 1 AOI31D1BWP7T $T=193040 82720 1 180 $X=188830 $Y=82485
X1643 1122 1128 402 1124 1061 2 1 AOI31D1BWP7T $T=194160 90560 0 0 $X=193870 $Y=90325
X1644 474 505 1142 514 1198 2 1 AOI31D1BWP7T $T=279840 67040 0 180 $X=275630 $Y=62830
X1645 523 521 1226 1223 412 2 1 AOI31D1BWP7T $T=282080 51360 0 180 $X=277870 $Y=47150
X1646 827 1 46 47 818 45 2 ND4D0BWP7T $T=41280 59200 0 180 $X=37630 $Y=54990
X1647 824 1 50 827 825 814 2 ND4D0BWP7T $T=41280 67040 1 180 $X=37630 $Y=66805
X1648 60 1 823 806 47 842 2 ND4D0BWP7T $T=41840 98400 0 0 $X=41550 $Y=98165
X1649 61 1 826 820 818 70 2 ND4D0BWP7T $T=41840 106240 1 0 $X=41550 $Y=102030
X1650 824 1 16 71 843 845 2 ND4D0BWP7T $T=43520 82720 0 0 $X=43230 $Y=82485
X1651 824 1 87 863 100 869 2 ND4D0BWP7T $T=53600 98400 1 0 $X=53310 $Y=94190
X1652 834 1 16 878 125 123 2 ND4D0BWP7T $T=61440 90560 0 0 $X=61150 $Y=90325
X1653 824 1 127 872 882 880 2 ND4D0BWP7T $T=63120 98400 1 0 $X=62830 $Y=94190
X1654 830 1 834 66 125 139 2 ND4D0BWP7T $T=65920 82720 1 0 $X=65630 $Y=78510
X1655 883 1 813 38 137 888 2 ND4D0BWP7T $T=66480 90560 0 0 $X=66190 $Y=90325
X1656 835 1 143 811 66 889 2 ND4D0BWP7T $T=69280 82720 0 0 $X=68990 $Y=82485
X1657 154 1 875 882 901 156 2 ND4D0BWP7T $T=80480 98400 1 0 $X=80190 $Y=94190
X1658 183 1 195 209 205 930 2 ND4D0BWP7T $T=101200 59200 1 180 $X=97550 $Y=58965
X1659 928 1 218 181 937 224 2 ND4D0BWP7T $T=101760 74880 1 0 $X=101470 $Y=70670
X1660 183 1 926 232 921 227 2 ND4D0BWP7T $T=108480 98400 0 180 $X=104830 $Y=94190
X1661 952 1 207 953 241 243 2 ND4D0BWP7T $T=107920 90560 1 0 $X=107630 $Y=86350
X1662 926 1 246 961 964 962 2 ND4D0BWP7T $T=111840 67040 0 0 $X=111550 $Y=66805
X1663 984 1 937 923 262 976 2 ND4D0BWP7T $T=128640 74880 0 180 $X=124990 $Y=70670
X1664 212 1 979 981 977 916 2 ND4D0BWP7T $T=128640 82720 0 180 $X=124990 $Y=78510
X1665 974 1 970 975 196 268 2 ND4D0BWP7T $T=125280 106240 1 0 $X=124990 $Y=102030
X1666 995 1 248 937 272 988 2 ND4D0BWP7T $T=133680 67040 1 180 $X=130030 $Y=66805
X1667 282 1 939 996 279 287 2 ND4D0BWP7T $T=136480 98400 1 180 $X=132830 $Y=98165
X1668 282 1 269 978 971 1000 2 ND4D0BWP7T $T=134240 67040 1 0 $X=133950 $Y=62830
X1669 199 1 952 970 999 290 2 ND4D0BWP7T $T=134800 90560 0 0 $X=134510 $Y=90325
X1670 251 1 995 269 292 1002 2 ND4D0BWP7T $T=136480 74880 1 0 $X=136190 $Y=70670
X1671 282 1 1010 1009 288 298 2 ND4D0BWP7T $T=144320 106240 0 180 $X=140670 $Y=102030
X1672 952 1 1007 1018 315 311 2 ND4D0BWP7T $T=146000 90560 0 0 $X=145710 $Y=90325
X1673 318 1 1017 971 306 1026 2 ND4D0BWP7T $T=148240 74880 0 0 $X=147950 $Y=74645
X1674 949 1 232 970 1009 1023 2 ND4D0BWP7T $T=157200 98400 0 180 $X=153550 $Y=94190
X1675 351 1 348 1042 1036 1037 2 ND4D0BWP7T $T=174000 82720 0 180 $X=170350 $Y=78510
X1676 367 1 1069 1066 360 1070 2 ND4D0BWP7T $T=180160 67040 0 180 $X=176510 $Y=62830
X1677 1067 1 1054 1073 1075 370 2 ND4D0BWP7T $T=177920 90560 1 0 $X=177630 $Y=86350
X1678 1106 1 1040 1071 381 1085 2 ND4D0BWP7T $T=189680 90560 0 180 $X=186030 $Y=86350
X1679 1121 1 1124 1120 1115 1087 2 ND4D0BWP7T $T=195280 82720 0 180 $X=191630 $Y=78510
X1680 1040 1 1121 400 1105 1129 2 ND4D0BWP7T $T=191920 90560 1 0 $X=191630 $Y=86350
X1681 1133 1 1036 1131 1075 1125 2 ND4D0BWP7T $T=198640 98400 0 180 $X=194990 $Y=94190
X1682 409 1 1140 1142 1039 1144 2 ND4D0BWP7T $T=207040 67040 1 0 $X=206750 $Y=62830
X1683 1106 1 419 1139 394 1138 2 ND4D0BWP7T $T=210960 98400 0 180 $X=207310 $Y=94190
X1684 1150 1 422 421 418 1135 2 ND4D0BWP7T $T=212080 51360 0 180 $X=208430 $Y=47150
X1685 1036 1 1154 1139 1156 1153 2 ND4D0BWP7T $T=211520 90560 0 0 $X=211230 $Y=90325
X1686 1161 1 431 1079 410 1152 2 ND4D0BWP7T $T=217680 74880 0 180 $X=214030 $Y=70670
X1687 1096 1 443 1166 1115 1162 2 ND4D0BWP7T $T=222720 67040 1 180 $X=219070 $Y=66805
X1688 1171 1 470 1170 1140 464 2 ND4D0BWP7T $T=238400 51360 0 180 $X=234750 $Y=47150
X1689 1176 1 1124 1154 1158 1199 2 ND4D0BWP7T $T=237840 82720 0 0 $X=237550 $Y=82485
X1690 134 1 906 2 153 159 IND3D1BWP7T $T=87760 51360 1 180 $X=84110 $Y=51125
X1691 346 1039 1095 2 1 NR2D1P5BWP7T $T=173440 59200 1 180 $X=169230 $Y=58965
X1692 1116 1073 398 2 1 NR2D1P5BWP7T $T=193600 67040 0 180 $X=189390 $Y=62830
X1693 1038 1139 457 2 1 NR2D1P5BWP7T $T=247920 59200 0 0 $X=247630 $Y=58965
X1694 1194 1213 1233 2 1 NR2D1P5BWP7T $T=289920 74880 0 0 $X=289630 $Y=74645
X1695 598 594 1262 2 1 NR2D1P5BWP7T $T=355440 98400 0 180 $X=351230 $Y=94190
X1696 598 637 643 2 1 NR2D1P5BWP7T $T=395200 98400 1 180 $X=390990 $Y=98165
X1697 314 304 1001 2 1 306 OA21D0BWP7T $T=148800 59200 0 180 $X=145150 $Y=54990
X1698 835 2 93 857 88 853 1 INR4D0BWP7T $T=55280 67040 0 180 $X=50510 $Y=62830
X1699 87 2 116 862 879 883 1 INR4D0BWP7T $T=59200 82720 1 0 $X=58910 $Y=78510
X1700 920 2 960 249 252 967 1 INR4D0BWP7T $T=110160 98400 1 0 $X=109870 $Y=94190
X1701 1028 2 283 931 192 1022 1 INR4D0BWP7T $T=155520 90560 1 180 $X=150750 $Y=90325
X1702 1040 2 352 1049 1048 1054 1 INR4D0BWP7T $T=170640 90560 0 0 $X=170350 $Y=90325
X1703 437 2 417 1119 1168 440 1 INR4D0BWP7T $T=218240 106240 1 0 $X=217950 $Y=102030
X1704 446 2 444 1111 1119 1165 1 INR4D0BWP7T $T=224400 82720 0 180 $X=219630 $Y=78510
X1705 1207 2 480 1114 1065 1190 1 INR4D0BWP7T $T=253520 51360 1 180 $X=248750 $Y=51125
X1706 837 1 57 829 2 833 IND3D0BWP7T $T=43520 82720 1 180 $X=39870 $Y=82485
X1707 1038 1 350 353 2 1055 IND3D0BWP7T $T=171200 51360 1 0 $X=170910 $Y=47150
X1708 1038 1 350 353 2 1057 IND3D0BWP7T $T=171200 51360 0 0 $X=170910 $Y=51125
X1709 1038 1 350 361 2 1064 IND3D0BWP7T $T=175120 51360 1 0 $X=174830 $Y=47150
X1710 1077 1 360 378 2 1076 IND3D0BWP7T $T=182960 51360 0 0 $X=182670 $Y=51125
X1711 807 1 822 814 817 2 NR3D1BWP7T $T=26720 74880 1 0 $X=26430 $Y=70670
X1712 78 1 864 138 151 2 NR3D1BWP7T $T=68720 98400 0 0 $X=68430 $Y=98165
X1713 936 1 208 930 941 2 NR3D1BWP7T $T=97840 67040 1 0 $X=97550 $Y=62830
X1714 1047 1 1048 1041 1036 2 NR3D1BWP7T $T=175120 74880 0 180 $X=170350 $Y=70670
X1715 356 1 352 1053 1066 2 NR3D1BWP7T $T=174000 82720 1 0 $X=173710 $Y=78510
X1716 1049 1 1082 1091 1072 2 NR3D1BWP7T $T=185760 90560 1 180 $X=180990 $Y=90325
X1717 389 1 391 1077 1115 2 NR3D1BWP7T $T=188560 59200 1 0 $X=188270 $Y=54990
X1718 415 1 1136 1146 1124 2 NR3D1BWP7T $T=210400 74880 1 180 $X=205630 $Y=74645
X1719 358 1 1163 1164 1105 2 NR3D1BWP7T $T=219360 90560 1 180 $X=214590 $Y=90325
X1720 441 1 1052 1167 394 2 NR3D1BWP7T $T=222720 98400 0 180 $X=217950 $Y=94190
X1721 812 1 820 811 39 53 2 IND4D0BWP7T $T=27280 98400 1 0 $X=26990 $Y=94190
X1722 150 1 54 868 136 856 2 IND4D0BWP7T $T=72080 98400 0 180 $X=67870 $Y=94190
X1723 890 1 901 100 898 905 2 IND4D0BWP7T $T=88320 98400 0 180 $X=84110 $Y=94190
X1724 890 1 868 906 908 899 2 IND4D0BWP7T $T=91120 82720 1 180 $X=86910 $Y=82485
X1725 244 1 246 181 963 251 2 IND4D0BWP7T $T=111280 51360 0 0 $X=110990 $Y=51125
X1726 213 1 986 921 990 957 2 IND4D0BWP7T $T=126960 90560 0 0 $X=126670 $Y=90325
X1727 1015 1 975 251 344 949 2 IND4D0BWP7T $T=166720 98400 0 0 $X=166430 $Y=98165
X1728 1116 1 1059 406 1130 409 2 IND4D0BWP7T $T=193600 67040 0 0 $X=193310 $Y=66805
X1729 457 1 1098 351 1174 1150 2 IND4D0BWP7T $T=229440 59200 1 180 $X=225230 $Y=58965
X1730 1149 1 1176 437 451 1180 2 IND4D0BWP7T $T=225520 98400 0 0 $X=225230 $Y=98165
X1731 862 1 870 830 101 846 2 IND4D1BWP7T $T=55280 74880 0 0 $X=54990 $Y=74645
X1732 105 1 129 91 885 835 2 IND4D1BWP7T $T=63680 90560 1 0 $X=63390 $Y=86350
X1733 946 1 236 240 225 245 2 IND4D1BWP7T $T=107360 106240 1 0 $X=107070 $Y=102030
X1734 372 1 423 1147 1132 409 2 IND4D1BWP7T $T=212640 51360 1 180 $X=207870 $Y=51125
X1735 1145 1 450 1173 1053 1040 2 IND4D1BWP7T $T=228320 74880 1 180 $X=223550 $Y=74645
X1736 1172 1 1179 406 1091 1184 2 IND4D1BWP7T $T=227760 90560 1 0 $X=227470 $Y=86350
X1737 78 52 837 848 828 1 2 INR4D1BWP7T $T=50240 74880 1 180 $X=43230 $Y=74645
X1738 191 213 943 219 226 1 2 INR4D1BWP7T $T=100640 82720 1 0 $X=100350 $Y=78510
X1739 988 991 982 266 216 1 2 INR4D1BWP7T $T=130880 67040 0 180 $X=123870 $Y=62830
X1740 364 1055 372 1067 377 1 2 INR4D1BWP7T $T=178480 51360 1 0 $X=178190 $Y=47150
X1741 1093 1102 1087 1094 350 1 2 INR4D1BWP7T $T=188000 82720 0 180 $X=180990 $Y=78510
X1742 436 438 1137 1131 1154 1 2 INR4D1BWP7T $T=219920 98400 1 180 $X=212910 $Y=98165
X1743 427 433 1164 1159 445 1 2 INR4D1BWP7T $T=216000 51360 0 0 $X=215710 $Y=51125
X1744 40 807 818 2 1 INR2D2BWP7T $T=31200 59200 0 180 $X=26430 $Y=54990
X1745 1188 1177 1179 2 1 INR2D2BWP7T $T=237840 82720 1 180 $X=233070 $Y=82485
X1746 6 2 11 1 15 NR2XD1BWP7T $T=21680 67040 1 0 $X=21390 $Y=62830
X1747 7 2 807 1 12 NR2XD1BWP7T $T=21680 90560 1 0 $X=21390 $Y=86350
X1748 7 2 18 1 23 NR2XD1BWP7T $T=22800 82720 0 0 $X=22510 $Y=82485
X1749 312 2 192 1 308 NR2XD1BWP7T $T=149920 74880 0 180 $X=145710 $Y=70670
X1750 312 2 321 1 319 NR2XD1BWP7T $T=152720 59200 0 180 $X=148510 $Y=54990
X1751 317 2 983 1 312 NR2XD1BWP7T $T=154960 51360 1 180 $X=150750 $Y=51125
X1752 465 2 446 1 1181 NR2XD1BWP7T $T=237280 90560 1 180 $X=233070 $Y=90325
X1753 1145 2 1128 1 1065 NR2XD1BWP7T $T=241200 67040 1 180 $X=236990 $Y=66805
X1754 1215 2 403 1 1195 NR2XD1BWP7T $T=262480 90560 1 180 $X=258270 $Y=90325
X1755 1201 2 1181 1 1224 NR2XD1BWP7T $T=266960 90560 1 0 $X=266670 $Y=86350
X1756 507 2 1043 1 1224 NR2XD1BWP7T $T=274800 82720 1 180 $X=270590 $Y=82485
X1757 1215 2 1111 1 506 NR2XD1BWP7T $T=277600 74880 0 180 $X=273390 $Y=70670
X1758 1215 2 1177 1 507 NR2XD1BWP7T $T=277600 82720 0 180 $X=273390 $Y=78510
X1759 503 2 1038 1 527 NR2XD1BWP7T $T=289920 51360 1 0 $X=289630 $Y=47150
X1760 1192 2 1223 1 525 NR2XD1BWP7T $T=293840 67040 0 180 $X=289630 $Y=62830
X1761 1192 2 472 1 1232 NR2XD1BWP7T $T=291600 59200 0 0 $X=291310 $Y=58965
X1762 1191 2 458 1 1194 NR2XD1BWP7T $T=299440 59200 0 180 $X=295230 $Y=54990
X1763 1227 2 496 1 1225 NR2XD1BWP7T $T=298880 59200 0 0 $X=298590 $Y=58965
X1764 33 1 816 804 2 IND2D1BWP7T $T=28960 74880 1 180 $X=25870 $Y=74645
X1765 807 1 881 79 2 IND2D1BWP7T $T=60880 59200 0 0 $X=60590 $Y=58965
X1766 99 1 891 140 2 IND2D1BWP7T $T=73200 90560 0 180 $X=70110 $Y=86350
X1767 283 1 297 338 2 IND2D1BWP7T $T=163920 98400 0 0 $X=163630 $Y=98165
X1768 442 1 1185 1170 2 IND2D1BWP7T $T=237280 67040 1 180 $X=234190 $Y=66805
X1769 490 1 1338 685 2 IND2D1BWP7T $T=432160 98400 1 0 $X=431870 $Y=94190
X1770 415 495 411 1181 2 1 1222 OR4XD1BWP7T $T=265280 82720 1 0 $X=264990 $Y=78510
X1771 368 1070 1068 1062 357 1 2 AO211D2BWP7T $T=180160 98400 1 180 $X=174830 $Y=98165
X1772 279 1 241 312 2 314 1019 OAI211D0BWP7T $T=146560 67040 1 0 $X=146270 $Y=62830
X1773 1100 1 1097 1090 2 375 1044 OAI211D0BWP7T $T=188000 106240 0 180 $X=184350 $Y=102030
X1774 1328 1 1324 1326 2 609 1329 OAI211D0BWP7T $T=420400 90560 0 180 $X=416750 $Y=86350
X1775 5 1 804 22 815 17 2 OAI211D2BWP7T $T=21120 67040 0 0 $X=20830 $Y=66805
X1776 1008 1 979 336 281 314 2 OAI211D2BWP7T $T=171200 67040 0 180 $X=164750 $Y=62830
X1777 1220 1 409 501 1155 1225 2 OAI211D2BWP7T $T=269200 74880 0 0 $X=268910 $Y=74645
X1778 251 1 247 959 2 CKND2D0BWP7T $T=112960 74880 0 0 $X=112670 $Y=74645
X1779 180 303 1011 294 1 2 1021 AO211D0BWP7T $T=143200 51360 0 0 $X=142910 $Y=51125
X1780 185 303 1019 962 1 2 1025 AO211D0BWP7T $T=153840 67040 0 180 $X=149630 $Y=62830
X1781 1213 1193 358 1114 1 2 1197 AO211D0BWP7T $T=258000 82720 1 180 $X=253790 $Y=82485
X1782 493 483 1214 1199 1 2 1211 AO211D0BWP7T $T=263040 82720 0 180 $X=258830 $Y=78510
X1783 805 2 803 813 810 19 1 AOI211D2BWP7T $T=21120 90560 0 0 $X=20830 $Y=90325
X1784 1060 2 444 1176 1186 1194 1 AOI211D2BWP7T $T=235040 74880 0 0 $X=234750 $Y=74645
X1785 499 2 411 1224 1 NR2D3BWP7T $T=267520 90560 0 0 $X=267230 $Y=90325
X1786 911 218 1 2 228 AN2D1BWP7T $T=103440 106240 1 0 $X=103150 $Y=102030
X1787 984 1008 1 2 932 AN2D1BWP7T $T=143760 74880 0 180 $X=140670 $Y=70670
X1788 10 811 4 1 2 ND2D2BWP7T $T=23920 51360 1 0 $X=23630 $Y=47150
X1789 187 184 177 1 2 ND2D2BWP7T $T=95600 51360 0 180 $X=91390 $Y=47150
X1790 423 415 1160 1 2 ND2D2BWP7T $T=217120 59200 0 180 $X=212910 $Y=54990
X1791 1186 409 481 1 2 ND2D2BWP7T $T=260240 74880 0 0 $X=259950 $Y=74645
X1792 1223 404 494 1 2 ND2D2BWP7T $T=275920 67040 0 180 $X=271710 $Y=62830
X1793 1232 1215 1213 1 2 ND2D2BWP7T $T=281520 82720 0 180 $X=277310 $Y=78510
X1794 608 2 1334 1309 659 1 653 1336 AOI221D1BWP7T $T=423760 82720 0 0 $X=423470 $Y=82485
X1795 68 1 2 808 72 843 NR3D0BWP7T $T=44080 90560 0 0 $X=43790 $Y=90325
X1796 858 1 2 97 80 852 NR3D0BWP7T $T=54720 67040 1 180 $X=51630 $Y=66805
X1797 107 1 2 864 98 850 NR3D0BWP7T $T=56400 98400 1 180 $X=53310 $Y=98165
X1798 116 1 2 108 58 106 NR3D0BWP7T $T=60320 90560 1 180 $X=57230 $Y=90325
X1799 1051 1 2 1046 1043 1035 NR3D0BWP7T $T=174560 67040 1 180 $X=171470 $Y=66805
X1800 1099 1 2 1076 1093 1090 NR3D0BWP7T $T=187440 98400 1 180 $X=184350 $Y=98165
X1801 386 1 2 1103 383 1083 NR3D0BWP7T $T=189680 51360 0 180 $X=186590 $Y=47150
X1802 1148 1 2 1127 414 1081 NR3D0BWP7T $T=209280 90560 1 180 $X=206190 $Y=90325
X1803 119 811 126 851 2 1 ND3D2BWP7T $T=60320 51360 1 0 $X=60030 $Y=47150
X1804 1232 1194 527 1225 2 1 ND3D2BWP7T $T=306720 51360 1 180 $X=301390 $Y=51125
X1805 959 2 235 997 1 NR2D0BWP7T $T=135360 82720 1 180 $X=132830 $Y=82485
X1806 16 806 828 124 133 1 2 ND4D2BWP7T $T=63680 74880 1 0 $X=63390 $Y=70670
X1807 153 73 148 90 158 1 2 ND4D2BWP7T $T=80480 51360 1 0 $X=80190 $Y=47150
X1808 205 193 911 184 201 1 2 ND4D2BWP7T $T=98960 98400 1 180 $X=91390 $Y=98165
X1809 920 928 226 949 944 1 2 ND4D2BWP7T $T=100640 67040 0 0 $X=100350 $Y=66805
X1810 952 940 933 183 229 1 2 ND4D2BWP7T $T=109600 90560 1 180 $X=102030 $Y=90325
X1811 135 1 130 880 68 816 2 OAI31D2BWP7T $T=68720 98400 1 180 $X=61710 $Y=98165
X1812 165 1 173 88 908 871 2 OAI31D2BWP7T $T=86640 90560 0 0 $X=86350 $Y=90325
X1813 824 1 46 852 2 85 ND3D1BWP7T $T=46880 90560 0 0 $X=46590 $Y=90325
X1814 67 1 91 31 2 862 ND3D1BWP7T $T=50240 90560 0 0 $X=49950 $Y=90325
X1815 43 1 67 835 2 99 ND3D1BWP7T $T=50800 82720 0 0 $X=50510 $Y=82485
X1816 117 1 834 811 2 93 ND3D1BWP7T $T=65920 82720 0 0 $X=65630 $Y=82485
X1817 212 1 929 932 2 203 ND3D1BWP7T $T=100640 82720 0 180 $X=96990 $Y=78510
X1818 209 1 937 210 2 211 ND3D1BWP7T $T=101760 74880 0 180 $X=98110 $Y=70670
X1819 1022 1 971 241 2 276 ND3D1BWP7T $T=150480 90560 0 180 $X=146830 $Y=86350
X1820 1109 1 1120 1139 2 416 ND3D1BWP7T $T=205920 59200 0 0 $X=205630 $Y=58965
X1821 439 1 1158 1156 2 1093 ND3D1BWP7T $T=220480 90560 0 180 $X=216830 $Y=86350
X1822 1203 1 431 1184 2 1141 ND3D1BWP7T $T=251280 67040 1 180 $X=247630 $Y=66805
X1823 25 2 52 810 1 832 9 AOI211D1BWP7T $T=41280 90560 1 180 $X=37630 $Y=90325
X1824 58 2 808 49 1 826 19 AOI211D1BWP7T $T=41840 106240 0 180 $X=38190 $Y=102030
X1825 859 2 80 59 1 849 77 AOI211D1BWP7T $T=50800 74880 0 180 $X=47150 $Y=70670
X1826 959 2 942 1031 1 1033 333 AOI211D1BWP7T $T=153840 82720 1 0 $X=153550 $Y=78510
X1827 337 2 969 322 1 1034 998 AOI211D1BWP7T $T=165040 82720 0 0 $X=164750 $Y=82485
X1828 1196 2 442 455 1 1204 496 AOI211D1BWP7T $T=267520 59200 1 180 $X=263870 $Y=58965
X1829 1283 2 594 605 1 1287 612 AOI211D1BWP7T $T=363840 98400 0 0 $X=363550 $Y=98165
X1830 1291 2 1288 620 1 1290 612 AOI211D1BWP7T $T=376160 98400 1 0 $X=375870 $Y=94190
X1831 1327 2 637 1325 1 1324 612 AOI211D1BWP7T $T=409200 98400 0 180 $X=405550 $Y=94190
X1832 204 1 269 212 284 997 2 IND4D2BWP7T $T=142080 82720 0 180 $X=133390 $Y=78510
X1833 806 2 863 78 1 INR2D1BWP7T $T=56400 90560 0 180 $X=53310 $Y=86350
X1834 404 2 1207 436 1 INR2D1BWP7T $T=251280 67040 1 0 $X=250990 $Y=62830
X1835 628 636 624 1311 608 1 2 640 AO221D0BWP7T $T=390160 51360 0 0 $X=389870 $Y=51125
X1836 1285 668 610 671 608 1 2 1335 AO221D0BWP7T $T=421520 98400 0 0 $X=421230 $Y=98165
X1838 537 1247 539 1249 2 1 561 DFCND1BWP7T $T=306720 90560 1 0 $X=306430 $Y=86350
X1839 537 1267 539 1263 2 1 1259 DFCND1BWP7T $T=350400 67040 0 180 $X=337230 $Y=62830
X1840 537 1271 539 1266 2 1 580 DFCND1BWP7T $T=351520 82720 1 180 $X=338350 $Y=82485
X1841 537 1275 539 1274 2 1 1253 DFCND1BWP7T $T=364960 51360 1 180 $X=351790 $Y=51125
X1842 537 1295 539 631 2 1 1308 DFCND1BWP7T $T=375040 51360 1 0 $X=374750 $Y=47150
X1843 537 1305 539 619 2 1 1286 DFCND1BWP7T $T=389040 74880 1 180 $X=375870 $Y=74645
X1844 537 1312 539 1261 2 1 1320 DFCND1BWP7T $T=390720 74880 0 0 $X=390430 $Y=74645
X1845 537 1322 539 1319 2 1 663 DFCND1BWP7T $T=430480 106240 0 180 $X=417310 $Y=102030
X1846 1241 536 341 1 2 XNR2D2BWP7T $T=305040 74880 0 180 $X=298030 $Y=70670
X1847 642 1307 535 1 2 XNR2D2BWP7T $T=396880 74880 0 180 $X=389870 $Y=70670
X1848 118 1 2 110 821 870 102 AOI211XD0BWP7T $T=60880 59200 0 180 $X=57230 $Y=54990
X1849 109 1 2 864 63 899 51 AOI211XD0BWP7T $T=83280 82720 1 180 $X=79630 $Y=82485
X1850 167 1 2 903 69 907 63 AOI211XD0BWP7T $T=90000 67040 1 180 $X=86350 $Y=66805
X1851 945 1 2 204 214 1005 300 AOI211XD0BWP7T $T=140960 59200 0 0 $X=140670 $Y=58965
X1852 316 1 2 274 322 1016 220 AOI211XD0BWP7T $T=149920 82720 0 0 $X=149630 $Y=82485
X1853 1114 1 2 352 486 1202 1213 AOI211XD0BWP7T $T=252960 74880 0 0 $X=252670 $Y=74645
X1854 1297 1 2 1288 623 1303 612 AOI211XD0BWP7T $T=381760 98400 1 0 $X=381470 $Y=94190
X1855 537 1252 539 544 1343 1 2 DFCND2BWP7T $T=321280 82720 1 180 $X=306430 $Y=82485
X1856 537 1269 539 1264 1260 1 2 DFCND2BWP7T $T=364400 74880 1 180 $X=349550 $Y=74645
X1857 537 1306 539 618 615 1 2 DFCND2BWP7T $T=389600 59200 0 180 $X=374750 $Y=54990
X1858 537 1313 539 1318 1321 1 2 DFCND2BWP7T $T=391280 67040 0 0 $X=390990 $Y=66805
X1859 804 1 26 13 7 2 OAI21D2BWP7T $T=21120 82720 1 0 $X=20830 $Y=78510
X1860 806 1 25 20 12 2 OAI21D2BWP7T $T=21680 98400 0 0 $X=21390 $Y=98165
X1861 910 1 921 185 917 2 OAI21D2BWP7T $T=89440 67040 1 0 $X=89150 $Y=62830
X1862 1079 1 1145 503 1215 2 OAI21D2BWP7T $T=274800 67040 1 180 $X=269470 $Y=66805
X1863 1092 375 1 1088 2 371 1080 OAI22D1BWP7T $T=185760 82720 1 180 $X=181550 $Y=82485
X1864 1279 609 1 591 2 1283 1281 OAI22D1BWP7T $T=366640 90560 1 180 $X=362430 $Y=90325
X1865 617 609 1 586 2 1297 1296 OAI22D1BWP7T $T=377840 90560 0 0 $X=377550 $Y=90325
X1866 161 1 2 909 DEL1BWP7T $T=94480 98400 0 180 $X=88590 $Y=94190
X1867 664 666 1323 1332 608 1 2 669 AO221D1BWP7T $T=418720 74880 0 0 $X=418430 $Y=74645
X1868 537 1240 539 1237 2 1 1231 DFCND0BWP7T $T=307280 106240 0 180 $X=294110 $Y=102030
X1869 537 1236 539 1238 2 1 553 DFCND0BWP7T $T=299440 98400 0 0 $X=299150 $Y=98165
X1870 537 1244 539 1246 2 1 558 DFCND0BWP7T $T=304480 90560 0 0 $X=304190 $Y=90325
X1871 537 584 539 1344 2 1 1251 DFCND0BWP7T $T=344800 59200 0 180 $X=331630 $Y=54990
X1872 537 600 539 585 2 1 1270 DFCND0BWP7T $T=358240 98400 1 180 $X=345070 $Y=98165
X1873 537 1278 539 1276 2 1 1273 DFCND0BWP7T $T=365520 67040 1 180 $X=352350 $Y=66805
X1874 537 1302 539 1292 2 1 1284 DFCND0BWP7T $T=388480 67040 0 180 $X=375310 $Y=62830
X1875 534 531 533 517 530 1238 2 1235 1 OA222D0BWP7T $T=299440 98400 0 180 $X=292990 $Y=94190
X1876 1242 531 540 538 530 513 2 1239 1 OA222D0BWP7T $T=304480 74880 1 180 $X=298030 $Y=74645
X1877 554 531 540 1238 530 1246 2 1245 1 OA222D0BWP7T $T=311760 98400 0 180 $X=305310 $Y=94190
X1878 1254 531 540 557 530 538 2 552 1 OA222D0BWP7T $T=319040 106240 0 180 $X=312590 $Y=102030
X1879 564 531 540 1246 530 1249 2 1248 1 OA222D0BWP7T $T=319600 82720 0 180 $X=313150 $Y=78510
X1880 576 531 540 1261 530 1263 2 1265 1 OA222D0BWP7T $T=334720 74880 1 0 $X=334430 $Y=70670
X1881 1272 531 540 1263 530 583 2 1268 1 OA222D0BWP7T $T=347040 59200 1 180 $X=340590 $Y=58965
X1882 1289 531 540 1266 530 1292 2 1298 1 OA222D0BWP7T $T=375600 67040 0 0 $X=375310 $Y=66805
X1883 630 531 533 1292 530 619 2 1294 1 OA222D0BWP7T $T=383440 82720 0 180 $X=376990 $Y=78510
X1884 650 531 540 641 530 646 2 644 1 OA222D0BWP7T $T=401920 51360 1 180 $X=395470 $Y=51125
X1885 1323 531 540 1319 530 1261 2 1316 1 OA222D0BWP7T $T=406400 82720 0 180 $X=399950 $Y=78510
X1886 655 531 540 652 530 641 2 651 1 OA222D0BWP7T $T=407520 106240 0 180 $X=401070 $Y=102030
X1887 658 531 540 654 530 618 2 1304 1 OA222D0BWP7T $T=409200 51360 1 180 $X=402750 $Y=51125
X1888 822 2 839 1 868 51 809 AOI211XD1BWP7T $T=50240 82720 1 0 $X=49950 $Y=78510
X1889 1027 2 1002 1 335 332 185 AOI211XD1BWP7T $T=170640 74880 0 180 $X=163630 $Y=70670
X1890 342 2 983 1 315 917 332 AOI211XD1BWP7T $T=170640 90560 1 180 $X=163630 $Y=90325
X1891 529 532 1 2 INVD2P5BWP7T $T=293840 90560 0 0 $X=293550 $Y=90325
X1892 579 581 1 2 INVD2P5BWP7T $T=337520 106240 1 0 $X=337230 $Y=102030
X1893 727 740 1 2 INVD2P5BWP7T $T=465760 90560 0 0 $X=465470 $Y=90325
X1894 737 738 1 2 INVD2P5BWP7T $T=468000 98400 1 0 $X=467710 $Y=94190
X1895 743 749 1 2 INVD2P5BWP7T $T=469680 51360 1 0 $X=469390 $Y=47150
X1896 531 551 1 533 544 530 1249 2 1252 OAI222D2BWP7T $T=311760 74880 0 0 $X=311470 $Y=74645
X1897 531 589 1 533 1264 530 577 2 1269 OAI222D2BWP7T $T=344800 74880 1 180 $X=334430 $Y=74645
X1898 531 578 1 540 571 530 583 2 590 OAI222D2BWP7T $T=335280 51360 0 0 $X=334990 $Y=51125
X1899 531 592 1 533 1266 530 585 2 1271 OAI222D2BWP7T $T=349280 90560 0 180 $X=338910 $Y=86350
X1900 531 1277 1 533 599 530 1264 2 1278 OAI222D2BWP7T $T=360480 67040 0 180 $X=350110 $Y=62830
X1901 531 1285 1 540 1274 530 571 2 1275 OAI222D2BWP7T $T=363840 51360 0 180 $X=353470 $Y=47150
X1902 531 1309 1 540 631 530 622 2 1295 OAI222D2BWP7T $T=388480 59200 1 180 $X=378110 $Y=58965
X1903 531 657 1 540 1318 530 1274 2 1313 OAI222D2BWP7T $T=406400 59200 1 180 $X=396030 $Y=58965
X1904 531 656 1 540 1319 530 649 2 1322 OAI222D2BWP7T $T=408640 98400 1 180 $X=398270 $Y=98165
X1905 531 674 1 540 667 530 1318 2 662 OAI222D2BWP7T $T=427680 59200 1 180 $X=417310 $Y=58965
X1906 389 401 1125 1126 405 1 2 OAI31D0BWP7T $T=192480 98400 0 0 $X=192190 $Y=98165
X1907 515 685 707 2 1 CKAN2D2BWP7T $T=443360 51360 0 0 $X=443070 $Y=51125
X1908 1201 1191 358 1154 2 1 IAO21D2BWP7T $T=252960 90560 0 180 $X=247630 $Y=86350
X1909 3 16 809 1 2 ND2D1P5BWP7T $T=22800 59200 1 0 $X=22510 $Y=54990
X1910 333 336 300 1 2 ND2D1P5BWP7T $T=164480 51360 1 0 $X=164190 $Y=47150
X1911 493 1195 535 1 2 ND2D1P5BWP7T $T=296080 67040 0 0 $X=295790 $Y=66805
X1912 186 918 928 190 1 2 206 IIND4D1BWP7T $T=93360 90560 1 0 $X=93070 $Y=86350
X1913 1024 2 1 910 330 NR2XD2BWP7T $T=149360 51360 1 0 $X=149070 $Y=47150
X1914 1 2 ICV_23 $T=77120 90560 0 0 $X=76830 $Y=90325
X1915 1 2 ICV_23 $T=134240 106240 1 0 $X=133950 $Y=102030
X1916 1 2 ICV_23 $T=166160 98400 1 0 $X=165870 $Y=94190
X1917 1 2 ICV_23 $T=168400 74880 0 0 $X=168110 $Y=74645
X1918 1 2 ICV_23 $T=195280 90560 1 0 $X=194990 $Y=86350
X1919 1 2 ICV_23 $T=227760 67040 0 0 $X=227470 $Y=66805
X1920 1 2 ICV_23 $T=245120 90560 0 0 $X=244830 $Y=90325
X1921 1 2 ICV_23 $T=252400 98400 1 0 $X=252110 $Y=94190
X1922 1 2 ICV_23 $T=263040 106240 1 0 $X=262750 $Y=102030
X1923 1 2 ICV_23 $T=279280 98400 1 0 $X=278990 $Y=94190
X1924 1 2 ICV_23 $T=287120 90560 1 0 $X=286830 $Y=86350
X1925 1 2 ICV_23 $T=300000 67040 0 0 $X=299710 $Y=66805
X1926 1 2 ICV_23 $T=307840 59200 1 0 $X=307550 $Y=54990
X1927 1 2 ICV_23 $T=311200 74880 1 0 $X=310910 $Y=70670
X1928 1 2 ICV_23 $T=321280 82720 0 0 $X=320990 $Y=82485
X1929 1 2 ICV_23 $T=329120 106240 1 0 $X=328830 $Y=102030
X1930 1 2 ICV_23 $T=363280 59200 1 0 $X=362990 $Y=54990
X1931 1 2 ICV_23 $T=371120 51360 0 0 $X=370830 $Y=51125
X1932 1 2 ICV_23 $T=413120 90560 0 0 $X=412830 $Y=90325
X1933 1 2 ICV_23 $T=427680 59200 0 0 $X=427390 $Y=58965
X1934 1 2 ICV_23 $T=447280 51360 0 0 $X=446990 $Y=51125
X1935 1 2 ICV_23 $T=447280 98400 1 0 $X=446990 $Y=94190
X1936 1 2 ICV_23 $T=455120 51360 0 0 $X=454830 $Y=51125
X1937 1 2 ICV_23 $T=455120 74880 1 0 $X=454830 $Y=70670
X1938 1 2 ICV_23 $T=461280 98400 1 0 $X=460990 $Y=94190
X1939 526 2 531 1 CKND10BWP7T $T=292160 82720 1 0 $X=291870 $Y=78510
X1940 597 606 1272 1256 608 611 1 2 AO221D2BWP7T $T=360480 59200 0 0 $X=360190 $Y=58965
X1941 614 634 1289 1314 608 648 1 2 AO221D2BWP7T $T=392400 90560 1 0 $X=392110 $Y=86350
X1942 1317 1 609 645 1315 586 2 OAI22D2BWP7T $T=402480 98400 0 180 $X=395470 $Y=94190
X1943 1088 1104 1101 1061 1094 2 1 OAI22D0BWP7T $T=189680 90560 1 180 $X=186030 $Y=90325
X1944 698 685 702 1 2 AN2D2BWP7T $T=442240 67040 0 0 $X=441950 $Y=66805
X1945 608 2 1277 1 679 NR2XD3BWP7T $T=432160 82720 0 180 $X=423470 $Y=78510
X1946 608 2 675 1 684 NR2XD3BWP7T $T=435520 74880 1 180 $X=426830 $Y=74645
X1947 608 2 1254 1 688 NR2XD3BWP7T $T=438880 90560 0 180 $X=430190 $Y=86350
X1948 608 2 687 1 705 NR2XD3BWP7T $T=444480 59200 1 180 $X=435790 $Y=58965
X1949 608 2 690 1 703 NR2XD3BWP7T $T=446720 74880 0 180 $X=438030 $Y=70670
X1950 608 2 678 1 701 NR2XD3BWP7T $T=446720 82720 0 180 $X=438030 $Y=78510
X1951 608 2 691 1 706 NR2XD3BWP7T $T=447280 82720 1 180 $X=438590 $Y=82485
X1952 608 2 692 1 704 NR2XD3BWP7T $T=447280 98400 0 180 $X=438590 $Y=94190
X1953 608 2 658 1 712 NR2XD3BWP7T $T=447840 59200 0 180 $X=439150 $Y=54990
X1954 608 2 694 1 715 NR2XD3BWP7T $T=448400 90560 1 180 $X=439710 $Y=90325
X1955 676 2 696 1 713 NR2XD3BWP7T $T=449520 74880 1 180 $X=440830 $Y=74645
X1956 676 2 697 1 710 NR2XD3BWP7T $T=450080 51360 0 180 $X=441390 $Y=47150
X1957 608 2 699 1 711 NR2XD3BWP7T $T=450080 90560 0 180 $X=441390 $Y=86350
X1958 676 2 721 1 742 NR2XD3BWP7T $T=468560 59200 1 180 $X=459870 $Y=58965
X1959 676 2 729 1 744 NR2XD3BWP7T $T=471920 74880 0 180 $X=463230 $Y=70670
X1960 676 2 731 1 747 NR2XD3BWP7T $T=472480 67040 0 180 $X=463790 $Y=62830
X1961 167 1 825 868 904 2 110 IIND4D0BWP7T $T=87760 67040 0 180 $X=82430 $Y=62830
X1962 1020 297 1010 999 2 977 1 IINR4D1BWP7T $T=151040 98400 1 180 $X=143470 $Y=98165
X1963 676 2 670 1 673 NR2D5BWP7T $T=431600 67040 0 180 $X=422910 $Y=62830
X1964 608 2 695 1 700 NR2D5BWP7T $T=448960 67040 0 180 $X=440270 $Y=62830
X1965 676 2 1242 1 723 NR2D5BWP7T $T=466880 67040 1 180 $X=458190 $Y=66805
X1966 676 672 665 1 2 INR2XD4BWP7T $T=432160 59200 0 180 $X=418990 $Y=54990
X1967 676 677 635 1 2 INR2XD4BWP7T $T=436080 51360 1 180 $X=422910 $Y=51125
X1968 676 683 642 1 2 INR2XD4BWP7T $T=440000 51360 0 180 $X=426830 $Y=47150
X1969 676 735 724 1 2 INR2XD4BWP7T $T=474160 59200 0 180 $X=460990 $Y=54990
X1970 257 1 960 2 972 OR2D1BWP7T $T=121920 90560 0 0 $X=121630 $Y=90325
X1971 1181 1 438 2 1049 OR2D1BWP7T $T=228320 90560 1 180 $X=225230 $Y=90325
X1972 453 1 452 2 1119 OR2D1BWP7T $T=228320 106240 0 180 $X=225230 $Y=102030
X1973 1198 1 393 2 466 OR2D1BWP7T $T=241200 106240 0 180 $X=238110 $Y=102030
X1974 1227 1 1191 2 1234 OR2D1BWP7T $T=279840 74880 0 0 $X=279550 $Y=74645
X1975 682 1 608 2 1337 OR2D1BWP7T $T=431040 106240 1 0 $X=430750 $Y=102030
X1976 689 1 608 2 1340 OR2D1BWP7T $T=438320 98400 0 0 $X=438030 $Y=98165
X1977 693 1 608 2 1341 OR2D1BWP7T $T=440000 106240 1 0 $X=439710 $Y=102030
X1978 1 2 ICV_33 $T=31200 59200 1 0 $X=30910 $Y=54990
X1979 1 2 ICV_33 $T=31200 67040 1 0 $X=30910 $Y=62830
X1980 1 2 ICV_33 $T=73200 98400 0 0 $X=72910 $Y=98165
X1981 1 2 ICV_33 $T=115200 59200 0 0 $X=114910 $Y=58965
X1982 1 2 ICV_33 $T=115200 82720 1 0 $X=114910 $Y=78510
X1983 1 2 ICV_33 $T=157200 59200 1 0 $X=156910 $Y=54990
X1984 1 2 ICV_33 $T=157200 59200 0 0 $X=156910 $Y=58965
X1985 1 2 ICV_33 $T=157200 67040 0 0 $X=156910 $Y=66805
X1986 1 2 ICV_33 $T=157200 82720 1 0 $X=156910 $Y=78510
X1987 1 2 ICV_33 $T=157200 82720 0 0 $X=156910 $Y=82485
X1988 1 2 ICV_33 $T=283200 90560 1 0 $X=282910 $Y=86350
X1989 1 2 ICV_33 $T=325200 82720 1 0 $X=324910 $Y=78510
X1990 1 2 ICV_33 $T=367200 90560 1 0 $X=366910 $Y=86350
X1991 1 2 ICV_33 $T=367200 98400 0 0 $X=366910 $Y=98165
X1992 1 2 ICV_33 $T=451200 74880 1 0 $X=450910 $Y=70670
X1993 1 2 ICV_33 $T=471360 67040 0 0 $X=471070 $Y=66805
X1994 1 2 ICV_34 $T=31200 74880 1 0 $X=30910 $Y=70670
X1995 1 2 ICV_34 $T=73200 59200 1 0 $X=72910 $Y=54990
X1996 1 2 ICV_34 $T=73200 59200 0 0 $X=72910 $Y=58965
X1997 1 2 ICV_34 $T=73200 67040 0 0 $X=72910 $Y=66805
X1998 1 2 ICV_34 $T=73200 90560 1 0 $X=72910 $Y=86350
X1999 1 2 ICV_34 $T=115200 67040 0 0 $X=114910 $Y=66805
X2000 1 2 ICV_34 $T=157200 74880 1 0 $X=156910 $Y=70670
X2001 1 2 ICV_34 $T=157200 98400 1 0 $X=156910 $Y=94190
X2002 1 2 ICV_34 $T=157200 106240 1 0 $X=156910 $Y=102030
X2003 1 2 ICV_34 $T=199200 98400 0 0 $X=198910 $Y=98165
X2004 1 2 ICV_34 $T=241200 59200 0 0 $X=240910 $Y=58965
X2005 1 2 ICV_34 $T=241200 74880 1 0 $X=240910 $Y=70670
X2006 1 2 ICV_34 $T=241200 90560 1 0 $X=240910 $Y=86350
X2007 1 2 ICV_34 $T=283200 67040 1 0 $X=282910 $Y=62830
X2008 1 2 ICV_34 $T=325200 67040 1 0 $X=324910 $Y=62830
X2009 1 2 ICV_34 $T=367200 98400 1 0 $X=366910 $Y=94190
X2010 1 2 ICV_34 $T=409200 98400 1 0 $X=408910 $Y=94190
X2011 1 2 ICV_34 $T=451200 82720 1 0 $X=450910 $Y=78510
.ENDS
***************************************
.SUBCKT ICV_36 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300 301
+ 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321
+ 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341
+ 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361
+ 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381
+ 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398
** N=549 EP=397 IP=3119 FDC=4438
M0 1 470 458 1 N L=1.8e-07 W=1e-06 $X=168075 $Y=28185 $D=0
M1 470 177 1 1 N L=1.8e-07 W=5e-07 $X=168880 $Y=28185 $D=0
M2 1 469 470 1 N L=1.8e-07 W=5e-07 $X=169600 $Y=28185 $D=0
M3 470 172 1 1 N L=1.8e-07 W=5e-07 $X=170400 $Y=28185 $D=0
M4 2 470 458 2 P L=1.8e-07 W=1.37e-06 $X=168400 $Y=30045 $D=16
M5 548 177 2 2 P L=1.8e-07 W=1.37e-06 $X=169200 $Y=30045 $D=16
M6 549 469 548 2 P L=1.8e-07 W=1.37e-06 $X=169800 $Y=30045 $D=16
M7 470 172 549 2 P L=1.8e-07 W=1.37e-06 $X=170400 $Y=30045 $D=16
X127 457 1 2 120 CKBD1BWP7T $T=102880 35680 0 0 $X=102590 $Y=35445
X128 508 1 2 264 CKBD1BWP7T $T=250720 35680 0 180 $X=248190 $Y=31470
X129 513 1 2 478 CKBD1BWP7T $T=280400 20000 1 180 $X=277870 $Y=19765
X130 355 1 2 542 CKBD1BWP7T $T=415920 27840 0 0 $X=415630 $Y=27605
X131 6 1 2 408 INVD0BWP7T $T=25600 27840 0 180 $X=23630 $Y=23630
X132 414 1 2 413 INVD0BWP7T $T=39600 27840 1 180 $X=37630 $Y=27605
X133 16 1 2 419 INVD0BWP7T $T=45760 27840 1 0 $X=45470 $Y=23630
X134 47 1 2 421 INVD0BWP7T $T=48560 27840 0 0 $X=48270 $Y=27605
X135 49 1 2 423 INVD0BWP7T $T=50240 35680 0 0 $X=49950 $Y=35445
X136 67 1 2 37 INVD0BWP7T $T=62000 43520 0 180 $X=60030 $Y=39310
X137 75 1 2 433 INVD0BWP7T $T=69280 43520 0 180 $X=67310 $Y=39310
X138 43 1 2 440 INVD0BWP7T $T=79920 35680 0 0 $X=79630 $Y=35445
X139 434 1 2 92 INVD0BWP7T $T=84400 27840 0 0 $X=84110 $Y=27605
X140 445 1 2 100 INVD0BWP7T $T=91680 43520 1 0 $X=91390 $Y=39310
X141 448 1 2 103 INVD0BWP7T $T=92240 43520 0 0 $X=91950 $Y=43285
X142 122 1 2 456 INVD0BWP7T $T=105680 20000 0 0 $X=105390 $Y=19765
X143 459 1 2 154 INVD0BWP7T $T=130880 43520 0 0 $X=130590 $Y=43285
X144 107 1 2 464 INVD0BWP7T $T=137040 35680 0 180 $X=135070 $Y=31470
X145 462 1 2 166 INVD0BWP7T $T=147120 43520 1 0 $X=146830 $Y=39310
X146 178 1 2 469 INVD0BWP7T $T=172320 35680 0 180 $X=170350 $Y=31470
X147 480 1 2 186 INVD0BWP7T $T=180160 35680 0 180 $X=178190 $Y=31470
X148 477 1 2 487 INVD0BWP7T $T=194160 35680 0 180 $X=192190 $Y=31470
X149 492 1 2 477 INVD0BWP7T $T=207600 35680 0 180 $X=205630 $Y=31470
X150 232 1 2 493 INVD0BWP7T $T=216000 35680 0 180 $X=214030 $Y=31470
X151 243 1 2 494 INVD0BWP7T $T=224400 43520 0 0 $X=224110 $Y=43285
X152 503 1 2 499 INVD0BWP7T $T=228320 27840 1 180 $X=226350 $Y=27605
X153 233 1 2 274 INVD0BWP7T $T=261920 43520 0 180 $X=259950 $Y=39310
X154 508 1 2 278 INVD0BWP7T $T=260800 35680 1 0 $X=260510 $Y=31470
X155 281 1 2 517 INVD0BWP7T $T=312880 43520 0 0 $X=312590 $Y=43285
X156 339 1 2 525 INVD0BWP7T $T=367200 43520 0 180 $X=365230 $Y=39310
X157 346 1 2 539 INVD0BWP7T $T=386240 35680 1 0 $X=385950 $Y=31470
X158 540 1 2 541 INVD0BWP7T $T=404720 35680 1 180 $X=402750 $Y=35445
X159 527 335 1 2 BUFFD1P5BWP7T $T=361040 35680 0 180 $X=357950 $Y=31470
X160 528 351 1 2 BUFFD1P5BWP7T $T=400800 27840 1 0 $X=400510 $Y=23630
X161 74 1 2 25 INVD3BWP7T $T=65920 20000 0 0 $X=65630 $Y=19765
X162 306 1 2 310 INVD3BWP7T $T=316800 35680 1 0 $X=316510 $Y=31470
X163 311 1 2 313 INVD3BWP7T $T=320720 35680 0 0 $X=320430 $Y=35445
X164 349 1 2 352 INVD3BWP7T $T=401920 35680 1 0 $X=401630 $Y=31470
X209 412 1 2 18 BUFFD1BWP7T $T=28960 27840 0 0 $X=28670 $Y=27605
X210 426 1 2 442 BUFFD1BWP7T $T=82160 27840 0 0 $X=81870 $Y=27605
X211 455 1 2 446 BUFFD1BWP7T $T=101760 20000 1 180 $X=99230 $Y=19765
X212 472 1 2 471 BUFFD1BWP7T $T=175120 27840 0 180 $X=172590 $Y=23630
X213 183 1 2 179 BUFFD1BWP7T $T=175680 43520 1 180 $X=173150 $Y=43285
X214 303 1 2 518 BUFFD1BWP7T $T=312320 35680 1 0 $X=312030 $Y=31470
X215 304 1 2 519 BUFFD1BWP7T $T=312880 27840 0 0 $X=312590 $Y=27605
X216 331 1 2 522 BUFFD1BWP7T $T=350960 27840 1 180 $X=348430 $Y=27605
X217 363 1 2 544 BUFFD1BWP7T $T=430480 35680 0 0 $X=430190 $Y=35445
X218 1 2 DCAP4BWP7T $T=58080 27840 1 0 $X=57790 $Y=23630
X219 1 2 DCAP4BWP7T $T=101760 43520 1 0 $X=101470 $Y=39310
X220 1 2 DCAP4BWP7T $T=132560 35680 0 0 $X=132270 $Y=35445
X221 1 2 DCAP4BWP7T $T=144880 43520 1 0 $X=144590 $Y=39310
X222 1 2 DCAP4BWP7T $T=153280 35680 1 0 $X=152990 $Y=31470
X223 1 2 DCAP4BWP7T $T=157760 20000 0 0 $X=157470 $Y=19765
X224 1 2 DCAP4BWP7T $T=171200 27840 0 0 $X=170910 $Y=27605
X225 1 2 DCAP4BWP7T $T=212080 27840 1 0 $X=211790 $Y=23630
X226 1 2 DCAP4BWP7T $T=226640 35680 1 0 $X=226350 $Y=31470
X227 1 2 DCAP4BWP7T $T=258560 35680 1 0 $X=258270 $Y=31470
X228 1 2 DCAP4BWP7T $T=261360 35680 0 0 $X=261070 $Y=35445
X229 1 2 DCAP4BWP7T $T=266960 35680 1 0 $X=266670 $Y=31470
X230 1 2 DCAP4BWP7T $T=275360 27840 0 0 $X=275070 $Y=27605
X231 1 2 DCAP4BWP7T $T=398560 27840 1 0 $X=398270 $Y=23630
X232 1 2 DCAP4BWP7T $T=409760 35680 1 0 $X=409470 $Y=31470
X233 1 2 DCAP4BWP7T $T=451760 35680 0 0 $X=451470 $Y=35445
X234 1 2 DCAP4BWP7T $T=459600 27840 1 0 $X=459310 $Y=23630
X235 1 2 DCAP4BWP7T $T=459600 35680 0 0 $X=459310 $Y=35445
X236 1 2 DCAP4BWP7T $T=468560 27840 1 0 $X=468270 $Y=23630
X237 1 2 ICV_3 $T=21120 27840 1 0 $X=20830 $Y=23630
X238 1 2 ICV_3 $T=24480 20000 0 0 $X=24190 $Y=19765
X239 1 2 ICV_3 $T=31200 27840 0 0 $X=30910 $Y=27605
X240 1 2 ICV_3 $T=31200 35680 1 0 $X=30910 $Y=31470
X241 1 2 ICV_3 $T=31200 35680 0 0 $X=30910 $Y=35445
X242 1 2 ICV_3 $T=31200 43520 0 0 $X=30910 $Y=43285
X243 1 2 ICV_3 $T=35120 20000 0 0 $X=34830 $Y=19765
X244 1 2 ICV_3 $T=35120 27840 0 0 $X=34830 $Y=27605
X245 1 2 ICV_3 $T=35120 35680 0 0 $X=34830 $Y=35445
X246 1 2 ICV_3 $T=35120 43520 1 0 $X=34830 $Y=39310
X247 1 2 ICV_3 $T=35120 43520 0 0 $X=34830 $Y=43285
X248 1 2 ICV_3 $T=57520 43520 1 0 $X=57230 $Y=39310
X249 1 2 ICV_3 $T=63120 20000 0 0 $X=62830 $Y=19765
X250 1 2 ICV_3 $T=73200 20000 0 0 $X=72910 $Y=19765
X251 1 2 ICV_3 $T=73200 43520 1 0 $X=72910 $Y=39310
X252 1 2 ICV_3 $T=77120 35680 1 0 $X=76830 $Y=31470
X253 1 2 ICV_3 $T=77120 43520 0 0 $X=76830 $Y=43285
X254 1 2 ICV_3 $T=115200 20000 0 0 $X=114910 $Y=19765
X255 1 2 ICV_3 $T=115200 43520 1 0 $X=114910 $Y=39310
X256 1 2 ICV_3 $T=119120 35680 1 0 $X=118830 $Y=31470
X257 1 2 ICV_3 $T=119120 43520 1 0 $X=118830 $Y=39310
X258 1 2 ICV_3 $T=144880 27840 0 0 $X=144590 $Y=27605
X259 1 2 ICV_3 $T=145440 35680 1 0 $X=145150 $Y=31470
X260 1 2 ICV_3 $T=157200 35680 1 0 $X=156910 $Y=31470
X261 1 2 ICV_3 $T=161120 35680 1 0 $X=160830 $Y=31470
X262 1 2 ICV_3 $T=179040 27840 0 0 $X=178750 $Y=27605
X263 1 2 ICV_3 $T=190800 43520 0 0 $X=190510 $Y=43285
X264 1 2 ICV_3 $T=192480 27840 1 0 $X=192190 $Y=23630
X265 1 2 ICV_3 $T=199200 35680 0 0 $X=198910 $Y=35445
X266 1 2 ICV_3 $T=203120 27840 0 0 $X=202830 $Y=27605
X267 1 2 ICV_3 $T=203120 35680 0 0 $X=202830 $Y=35445
X268 1 2 ICV_3 $T=212640 35680 0 0 $X=212350 $Y=35445
X269 1 2 ICV_3 $T=222720 43520 1 0 $X=222430 $Y=39310
X270 1 2 ICV_3 $T=230000 43520 1 0 $X=229710 $Y=39310
X271 1 2 ICV_3 $T=230560 27840 0 0 $X=230270 $Y=27605
X272 1 2 ICV_3 $T=256880 27840 1 0 $X=256590 $Y=23630
X273 1 2 ICV_3 $T=287120 35680 1 0 $X=286830 $Y=31470
X274 1 2 ICV_3 $T=298320 20000 0 0 $X=298030 $Y=19765
X275 1 2 ICV_3 $T=312320 27840 1 0 $X=312030 $Y=23630
X276 1 2 ICV_3 $T=333600 27840 0 0 $X=333310 $Y=27605
X277 1 2 ICV_3 $T=357120 27840 1 0 $X=356830 $Y=23630
X278 1 2 ICV_3 $T=371120 27840 0 0 $X=370830 $Y=27605
X279 1 2 ICV_3 $T=409200 20000 0 0 $X=408910 $Y=19765
X280 1 2 ICV_3 $T=409200 35680 0 0 $X=408910 $Y=35445
X281 1 2 ICV_3 $T=413120 20000 0 0 $X=412830 $Y=19765
X282 1 2 ICV_3 $T=413120 27840 0 0 $X=412830 $Y=27605
X283 1 2 ICV_3 $T=432720 20000 0 0 $X=432430 $Y=19765
X284 1 2 ICV_3 $T=444480 27840 0 0 $X=444190 $Y=27605
X285 1 2 ICV_3 $T=459600 20000 0 0 $X=459310 $Y=19765
X286 1 2 DCAP8BWP7T $T=23360 43520 0 0 $X=23070 $Y=43285
X287 1 2 DCAP8BWP7T $T=29520 27840 1 0 $X=29230 $Y=23630
X288 1 2 DCAP8BWP7T $T=70400 35680 1 0 $X=70110 $Y=31470
X289 1 2 DCAP8BWP7T $T=70400 35680 0 0 $X=70110 $Y=35445
X290 1 2 DCAP8BWP7T $T=77120 27840 0 0 $X=76830 $Y=27605
X291 1 2 DCAP8BWP7T $T=94480 27840 1 0 $X=94190 $Y=23630
X292 1 2 DCAP8BWP7T $T=103440 27840 1 0 $X=103150 $Y=23630
X293 1 2 DCAP8BWP7T $T=112960 27840 1 0 $X=112670 $Y=23630
X294 1 2 DCAP8BWP7T $T=119120 27840 1 0 $X=118830 $Y=23630
X295 1 2 DCAP8BWP7T $T=119120 43520 0 0 $X=118830 $Y=43285
X296 1 2 DCAP8BWP7T $T=128080 20000 0 0 $X=127790 $Y=19765
X297 1 2 DCAP8BWP7T $T=137040 35680 1 0 $X=136750 $Y=31470
X298 1 2 DCAP8BWP7T $T=147680 35680 0 0 $X=147390 $Y=35445
X299 1 2 DCAP8BWP7T $T=153280 20000 0 0 $X=152990 $Y=19765
X300 1 2 DCAP8BWP7T $T=153840 43520 1 0 $X=153550 $Y=39310
X301 1 2 DCAP8BWP7T $T=166160 35680 1 0 $X=165870 $Y=31470
X302 1 2 DCAP8BWP7T $T=167280 20000 0 0 $X=166990 $Y=19765
X303 1 2 DCAP8BWP7T $T=168400 27840 1 0 $X=168110 $Y=23630
X304 1 2 DCAP8BWP7T $T=175120 27840 1 0 $X=174830 $Y=23630
X305 1 2 DCAP8BWP7T $T=175680 43520 0 0 $X=175390 $Y=43285
X306 1 2 DCAP8BWP7T $T=186320 43520 0 0 $X=186030 $Y=43285
X307 1 2 DCAP8BWP7T $T=188560 35680 0 0 $X=188270 $Y=35445
X308 1 2 DCAP8BWP7T $T=194160 35680 1 0 $X=193870 $Y=31470
X309 1 2 DCAP8BWP7T $T=196400 43520 1 0 $X=196110 $Y=39310
X310 1 2 DCAP8BWP7T $T=217680 27840 1 0 $X=217390 $Y=23630
X311 1 2 DCAP8BWP7T $T=239520 35680 1 0 $X=239230 $Y=31470
X312 1 2 DCAP8BWP7T $T=245120 43520 0 0 $X=244830 $Y=43285
X313 1 2 DCAP8BWP7T $T=262480 35680 1 0 $X=262190 $Y=31470
X314 1 2 DCAP8BWP7T $T=279840 35680 0 0 $X=279550 $Y=35445
X315 1 2 DCAP8BWP7T $T=280400 20000 0 0 $X=280110 $Y=19765
X316 1 2 DCAP8BWP7T $T=280960 43520 0 0 $X=280670 $Y=43285
X317 1 2 DCAP8BWP7T $T=281520 27840 0 0 $X=281230 $Y=27605
X318 1 2 DCAP8BWP7T $T=296080 27840 1 0 $X=295790 $Y=23630
X319 1 2 DCAP8BWP7T $T=302800 20000 0 0 $X=302510 $Y=19765
X320 1 2 DCAP8BWP7T $T=302800 35680 0 0 $X=302510 $Y=35445
X321 1 2 DCAP8BWP7T $T=307840 27840 1 0 $X=307550 $Y=23630
X322 1 2 DCAP8BWP7T $T=314560 43520 0 0 $X=314270 $Y=43285
X323 1 2 DCAP8BWP7T $T=342000 20000 0 0 $X=341710 $Y=19765
X324 1 2 DCAP8BWP7T $T=349280 20000 0 0 $X=348990 $Y=19765
X325 1 2 DCAP8BWP7T $T=349840 35680 1 0 $X=349550 $Y=31470
X326 1 2 DCAP8BWP7T $T=352640 27840 1 0 $X=352350 $Y=23630
X327 1 2 DCAP8BWP7T $T=362160 20000 0 0 $X=361870 $Y=19765
X328 1 2 DCAP8BWP7T $T=363840 35680 0 0 $X=363550 $Y=35445
X329 1 2 DCAP8BWP7T $T=384000 20000 0 0 $X=383710 $Y=19765
X330 1 2 DCAP8BWP7T $T=391840 43520 0 0 $X=391550 $Y=43285
X331 1 2 DCAP8BWP7T $T=396880 35680 1 0 $X=396590 $Y=31470
X332 1 2 DCAP8BWP7T $T=403600 27840 1 0 $X=403310 $Y=23630
X333 1 2 DCAP8BWP7T $T=404720 20000 0 0 $X=404430 $Y=19765
X334 1 2 DCAP8BWP7T $T=404720 35680 0 0 $X=404430 $Y=35445
X335 1 2 DCAP8BWP7T $T=405840 43520 0 0 $X=405550 $Y=43285
X336 1 2 DCAP8BWP7T $T=407520 43520 1 0 $X=407230 $Y=39310
X337 1 2 DCAP8BWP7T $T=422080 43520 1 0 $X=421790 $Y=39310
X338 1 2 DCAP8BWP7T $T=428240 20000 0 0 $X=427950 $Y=19765
X339 1 2 DCAP8BWP7T $T=440000 27840 0 0 $X=439710 $Y=27605
X340 1 2 DCAP8BWP7T $T=440560 43520 1 0 $X=440270 $Y=39310
X341 1 2 DCAP8BWP7T $T=441120 27840 1 0 $X=440830 $Y=23630
X342 1 2 DCAP8BWP7T $T=445600 20000 0 0 $X=445310 $Y=19765
X343 1 2 DCAP8BWP7T $T=447280 35680 0 0 $X=446990 $Y=35445
X344 1 2 DCAP8BWP7T $T=447840 35680 1 0 $X=447550 $Y=31470
X345 1 2 DCAP8BWP7T $T=448960 27840 1 0 $X=448670 $Y=23630
X346 1 2 DCAP8BWP7T $T=448960 43520 1 0 $X=448670 $Y=39310
X347 1 2 DCAP8BWP7T $T=449520 27840 0 0 $X=449230 $Y=27605
X348 1 2 DCAP8BWP7T $T=455120 27840 1 0 $X=454830 $Y=23630
X349 1 2 DCAP8BWP7T $T=460720 27840 0 0 $X=460430 $Y=27605
X350 1 2 DCAP8BWP7T $T=468000 35680 1 0 $X=467710 $Y=31470
X351 2 1 DCAPBWP7T $T=60320 27840 0 0 $X=60030 $Y=27605
X352 2 1 DCAPBWP7T $T=81600 20000 0 0 $X=81310 $Y=19765
X353 2 1 DCAPBWP7T $T=90000 35680 0 0 $X=89710 $Y=35445
X354 2 1 DCAPBWP7T $T=90560 43520 0 0 $X=90270 $Y=43285
X355 2 1 DCAPBWP7T $T=91680 27840 0 0 $X=91390 $Y=27605
X356 2 1 DCAPBWP7T $T=95040 27840 0 0 $X=94750 $Y=27605
X357 2 1 DCAPBWP7T $T=104560 27840 0 0 $X=104270 $Y=27605
X358 2 1 DCAPBWP7T $T=129200 27840 0 0 $X=128910 $Y=27605
X359 2 1 DCAPBWP7T $T=141520 35680 1 0 $X=141230 $Y=31470
X360 2 1 DCAPBWP7T $T=158320 43520 1 0 $X=158030 $Y=39310
X361 2 1 DCAPBWP7T $T=165600 27840 0 0 $X=165310 $Y=27605
X362 2 1 DCAPBWP7T $T=184080 27840 0 0 $X=183790 $Y=27605
X363 2 1 DCAPBWP7T $T=188560 27840 1 0 $X=188270 $Y=23630
X364 2 1 DCAPBWP7T $T=189120 43520 1 0 $X=188830 $Y=39310
X365 2 1 DCAPBWP7T $T=209840 43520 1 0 $X=209550 $Y=39310
X366 2 1 DCAPBWP7T $T=249600 43520 0 0 $X=249310 $Y=43285
X367 2 1 DCAPBWP7T $T=265840 43520 1 0 $X=265550 $Y=39310
X368 2 1 DCAPBWP7T $T=276480 20000 0 0 $X=276190 $Y=19765
X369 2 1 DCAPBWP7T $T=276480 35680 1 0 $X=276190 $Y=31470
X370 2 1 DCAPBWP7T $T=284320 35680 0 0 $X=284030 $Y=35445
X371 2 1 DCAPBWP7T $T=291600 20000 0 0 $X=291310 $Y=19765
X372 2 1 DCAPBWP7T $T=297200 35680 0 0 $X=296910 $Y=35445
X373 2 1 DCAPBWP7T $T=303360 43520 0 0 $X=303070 $Y=43285
X374 2 1 DCAPBWP7T $T=304480 43520 1 0 $X=304190 $Y=39310
X375 2 1 DCAPBWP7T $T=307280 20000 0 0 $X=306990 $Y=19765
X376 2 1 DCAPBWP7T $T=326320 35680 0 0 $X=326030 $Y=35445
X377 2 1 DCAPBWP7T $T=347040 27840 1 0 $X=346750 $Y=23630
X378 2 1 DCAPBWP7T $T=353760 20000 0 0 $X=353470 $Y=19765
X379 2 1 DCAPBWP7T $T=368320 35680 0 0 $X=368030 $Y=35445
X380 2 1 DCAPBWP7T $T=368320 43520 0 0 $X=368030 $Y=43285
X381 2 1 DCAPBWP7T $T=375600 20000 0 0 $X=375310 $Y=19765
X382 2 1 DCAPBWP7T $T=375600 35680 1 0 $X=375310 $Y=31470
X383 2 1 DCAPBWP7T $T=380080 43520 0 0 $X=379790 $Y=43285
X384 2 1 DCAPBWP7T $T=384560 35680 1 0 $X=384270 $Y=31470
X385 2 1 DCAPBWP7T $T=410320 43520 0 0 $X=410030 $Y=43285
X386 2 1 DCAPBWP7T $T=432720 35680 0 0 $X=432430 $Y=35445
X387 2 1 DCAPBWP7T $T=437200 27840 1 0 $X=436910 $Y=23630
X388 2 1 DCAPBWP7T $T=452320 35680 1 0 $X=452030 $Y=31470
X389 2 1 DCAPBWP7T $T=472480 35680 1 0 $X=472190 $Y=31470
X390 1 2 ICV_4 $T=41840 35680 1 0 $X=41550 $Y=31470
X391 1 2 ICV_4 $T=102880 43520 0 0 $X=102590 $Y=43285
X392 1 2 ICV_4 $T=119120 27840 0 0 $X=118830 $Y=27605
X393 1 2 ICV_4 $T=139840 20000 0 0 $X=139550 $Y=19765
X394 1 2 ICV_4 $T=156080 35680 0 0 $X=155790 $Y=35445
X395 1 2 ICV_4 $T=169520 43520 0 0 $X=169230 $Y=43285
X396 1 2 ICV_4 $T=268640 20000 0 0 $X=268350 $Y=19765
X397 1 2 ICV_4 $T=282080 35680 1 0 $X=281790 $Y=31470
X398 1 2 ICV_4 $T=282080 43520 1 0 $X=281790 $Y=39310
X399 1 2 ICV_4 $T=287120 35680 0 0 $X=286830 $Y=35445
X400 1 2 ICV_4 $T=287120 43520 1 0 $X=286830 $Y=39310
X401 1 2 ICV_4 $T=296640 43520 1 0 $X=296350 $Y=39310
X402 1 2 ICV_4 $T=299440 35680 1 0 $X=299150 $Y=31470
X403 1 2 ICV_4 $T=308400 35680 1 0 $X=308110 $Y=31470
X404 1 2 ICV_4 $T=324080 43520 1 0 $X=323790 $Y=39310
X405 1 2 ICV_4 $T=329120 43520 0 0 $X=328830 $Y=43285
X406 1 2 ICV_4 $T=333600 35680 1 0 $X=333310 $Y=31470
X407 1 2 ICV_4 $T=408080 27840 1 0 $X=407790 $Y=23630
X408 1 2 ICV_4 $T=408080 27840 0 0 $X=407790 $Y=27605
X409 1 2 ICV_4 $T=450080 20000 0 0 $X=449790 $Y=19765
X410 319 320 323 2 1 521 DFCNQD1BWP7T $T=333600 35680 0 0 $X=333310 $Y=35445
X411 319 325 323 2 1 523 DFCNQD1BWP7T $T=337520 35680 1 0 $X=337230 $Y=31470
X412 319 334 323 2 1 526 DFCNQD1BWP7T $T=353200 43520 1 0 $X=352910 $Y=39310
X413 319 359 323 2 1 528 DFCNQD1BWP7T $T=428240 20000 1 180 $X=415630 $Y=19765
X414 319 361 323 2 1 543 DFCNQD1BWP7T $T=429920 35680 0 180 $X=417310 $Y=31470
X535 1 2 ICV_9 $T=34000 35680 1 0 $X=33710 $Y=31470
X536 1 2 ICV_9 $T=76000 20000 0 0 $X=75710 $Y=19765
X537 1 2 ICV_9 $T=118000 20000 0 0 $X=117710 $Y=19765
X538 1 2 ICV_9 $T=160000 27840 0 0 $X=159710 $Y=27605
X539 1 2 ICV_9 $T=160000 35680 0 0 $X=159710 $Y=35445
X540 1 2 ICV_9 $T=286000 20000 0 0 $X=285710 $Y=19765
X541 1 2 ICV_9 $T=286000 27840 1 0 $X=285710 $Y=23630
X542 1 2 ICV_9 $T=286000 27840 0 0 $X=285710 $Y=27605
X543 1 2 ICV_9 $T=328000 20000 0 0 $X=327710 $Y=19765
X544 1 2 ICV_9 $T=328000 27840 0 0 $X=327710 $Y=27605
X545 1 2 ICV_9 $T=328000 35680 1 0 $X=327710 $Y=31470
X546 1 2 ICV_9 $T=328000 35680 0 0 $X=327710 $Y=35445
X547 1 2 ICV_9 $T=370000 20000 0 0 $X=369710 $Y=19765
X548 1 2 ICV_9 $T=370000 27840 1 0 $X=369710 $Y=23630
X549 1 2 ICV_9 $T=370000 35680 1 0 $X=369710 $Y=31470
X550 1 2 ICV_9 $T=412000 35680 1 0 $X=411710 $Y=31470
X551 1 2 ICV_9 $T=412000 35680 0 0 $X=411710 $Y=35445
X552 1 2 ICV_9 $T=454000 20000 0 0 $X=453710 $Y=19765
X553 1 2 ICV_9 $T=454000 35680 0 0 $X=453710 $Y=35445
X554 1 2 ICV_9 $T=454000 43520 0 0 $X=453710 $Y=43285
X574 1 2 ICV_13 $T=21120 43520 1 0 $X=20830 $Y=39310
X575 1 2 ICV_13 $T=30640 43520 1 0 $X=30350 $Y=39310
X576 1 2 ICV_13 $T=35120 27840 1 0 $X=34830 $Y=23630
X577 1 2 ICV_13 $T=42400 27840 1 0 $X=42110 $Y=23630
X578 1 2 ICV_13 $T=77120 43520 1 0 $X=76830 $Y=39310
X579 1 2 ICV_13 $T=87200 35680 1 0 $X=86910 $Y=31470
X580 1 2 ICV_13 $T=129200 27840 1 0 $X=128910 $Y=23630
X581 1 2 ICV_13 $T=156640 27840 1 0 $X=156350 $Y=23630
X582 1 2 ICV_13 $T=156640 27840 0 0 $X=156350 $Y=27605
X583 1 2 ICV_13 $T=156640 43520 0 0 $X=156350 $Y=43285
X584 1 2 ICV_13 $T=161120 20000 0 0 $X=160830 $Y=19765
X585 1 2 ICV_13 $T=161120 27840 1 0 $X=160830 $Y=23630
X586 1 2 ICV_13 $T=161120 43520 0 0 $X=160830 $Y=43285
X587 1 2 ICV_13 $T=172320 35680 1 0 $X=172030 $Y=31470
X588 1 2 ICV_13 $T=187440 27840 0 0 $X=187150 $Y=27605
X589 1 2 ICV_13 $T=198640 27840 1 0 $X=198350 $Y=23630
X590 1 2 ICV_13 $T=198640 35680 1 0 $X=198350 $Y=31470
X591 1 2 ICV_13 $T=215440 43520 1 0 $X=215150 $Y=39310
X592 1 2 ICV_13 $T=221040 43520 0 0 $X=220750 $Y=43285
X593 1 2 ICV_13 $T=222160 27840 1 0 $X=221870 $Y=23630
X594 1 2 ICV_13 $T=245120 20000 0 0 $X=244830 $Y=19765
X595 1 2 ICV_13 $T=245120 35680 1 0 $X=244830 $Y=31470
X596 1 2 ICV_13 $T=249600 27840 1 0 $X=249310 $Y=23630
X597 1 2 ICV_13 $T=256320 43520 1 0 $X=256030 $Y=39310
X598 1 2 ICV_13 $T=282640 27840 1 0 $X=282350 $Y=23630
X599 1 2 ICV_13 $T=300560 27840 1 0 $X=300270 $Y=23630
X600 1 2 ICV_13 $T=308960 43520 0 0 $X=308670 $Y=43285
X601 1 2 ICV_13 $T=324640 20000 0 0 $X=324350 $Y=19765
X602 1 2 ICV_13 $T=324640 35680 1 0 $X=324350 $Y=31470
X603 1 2 ICV_13 $T=324640 43520 0 0 $X=324350 $Y=43285
X604 1 2 ICV_13 $T=366640 20000 0 0 $X=366350 $Y=19765
X605 1 2 ICV_13 $T=366640 35680 1 0 $X=366350 $Y=31470
X606 1 2 ICV_13 $T=371120 43520 1 0 $X=370830 $Y=39310
X607 1 2 ICV_13 $T=388480 20000 0 0 $X=388190 $Y=19765
X608 1 2 ICV_13 $T=396320 43520 0 0 $X=396030 $Y=43285
X609 1 2 ICV_13 $T=413120 43520 0 0 $X=412830 $Y=43285
X610 1 2 ICV_13 $T=450640 43520 0 0 $X=450350 $Y=43285
X611 1 2 ICV_13 $T=455120 27840 0 0 $X=454830 $Y=27605
X612 1 2 ICV_13 $T=464080 43520 1 0 $X=463790 $Y=39310
X613 1 2 ICV_13 $T=465200 27840 0 0 $X=464910 $Y=27605
X614 1 2 ICV_13 $T=470800 27840 0 0 $X=470510 $Y=27605
X615 1 2 ICV_13 $T=470800 43520 0 0 $X=470510 $Y=43285
X616 410 1 2 19 INVD1BWP7T $T=29520 35680 0 0 $X=29230 $Y=35445
X617 39 1 2 416 INVD1BWP7T $T=45760 35680 1 0 $X=45470 $Y=31470
X618 28 1 2 12 INVD1BWP7T $T=50240 35680 1 180 $X=48270 $Y=35445
X619 45 1 2 24 INVD1BWP7T $T=58080 35680 0 0 $X=57790 $Y=35445
X620 46 1 2 65 INVD1BWP7T $T=58640 35680 1 0 $X=58350 $Y=31470
X621 431 1 2 81 INVD1BWP7T $T=81600 35680 1 0 $X=81310 $Y=31470
X622 409 1 2 87 INVD1BWP7T $T=83840 43520 1 180 $X=81870 $Y=43285
X623 52 1 2 437 INVD1BWP7T $T=86080 27840 0 0 $X=85790 $Y=27605
X624 101 1 2 105 INVD1BWP7T $T=93360 27840 0 0 $X=93070 $Y=27605
X625 108 1 2 447 INVD1BWP7T $T=99520 35680 0 180 $X=97550 $Y=31470
X626 110 1 2 112 INVD1BWP7T $T=101760 43520 0 180 $X=99790 $Y=39310
X627 453 1 2 452 INVD1BWP7T $T=100640 27840 0 0 $X=100350 $Y=27605
X628 139 1 2 451 INVD1BWP7T $T=110720 35680 0 180 $X=108750 $Y=31470
X629 137 1 2 449 INVD1BWP7T $T=115200 43520 0 180 $X=113230 $Y=39310
X630 138 1 2 133 INVD1BWP7T $T=115200 43520 1 180 $X=113230 $Y=43285
X631 466 1 2 461 INVD1BWP7T $T=143200 43520 0 180 $X=141230 $Y=39310
X632 145 1 2 157 INVD1BWP7T $T=144880 43520 0 180 $X=142910 $Y=39310
X633 467 1 2 465 INVD1BWP7T $T=143760 20000 0 0 $X=143470 $Y=19765
X634 164 1 2 143 INVD1BWP7T $T=147680 43520 1 180 $X=145710 $Y=43285
X635 156 1 2 173 INVD1BWP7T $T=157200 35680 0 180 $X=155230 $Y=31470
X636 475 1 2 187 INVD1BWP7T $T=175680 35680 1 0 $X=175390 $Y=31470
X637 193 1 2 191 INVD1BWP7T $T=181840 43520 0 180 $X=179870 $Y=39310
X638 260 1 2 236 INVD1BWP7T $T=232240 35680 1 180 $X=230270 $Y=35445
X639 246 1 2 251 INVD1BWP7T $T=232240 43520 1 180 $X=230270 $Y=43285
X640 509 1 2 484 INVD1BWP7T $T=250160 35680 1 180 $X=248190 $Y=35445
X641 270 1 2 242 INVD1BWP7T $T=254640 35680 0 180 $X=252670 $Y=31470
X642 276 1 2 505 INVD1BWP7T $T=261360 43520 1 180 $X=259390 $Y=43285
X643 280 1 2 262 INVD1BWP7T $T=265840 43520 0 180 $X=263870 $Y=39310
X644 272 1 2 286 INVD1BWP7T $T=270880 43520 0 0 $X=270590 $Y=43285
X645 252 1 2 511 INVD1BWP7T $T=293840 27840 1 180 $X=291870 $Y=27605
X646 514 1 2 479 INVD1BWP7T $T=296640 43520 0 180 $X=294670 $Y=39310
X647 294 1 2 291 INVD1BWP7T $T=302800 20000 1 180 $X=300830 $Y=19765
X648 298 1 2 516 INVD1BWP7T $T=311760 35680 1 180 $X=309790 $Y=35445
X649 525 1 2 524 INVD1BWP7T $T=356000 35680 0 180 $X=354030 $Y=31470
X650 524 1 2 529 INVD1BWP7T $T=373920 27840 0 0 $X=373630 $Y=27605
X651 351 1 2 356 INVD1BWP7T $T=418160 43520 1 180 $X=416190 $Y=43285
X652 521 322 1 2 BUFFD2BWP7T $T=339760 27840 1 180 $X=336110 $Y=27605
X653 526 314 1 2 BUFFD2BWP7T $T=356000 43520 0 0 $X=355710 $Y=43285
X654 543 357 1 2 BUFFD2BWP7T $T=417600 35680 0 0 $X=417310 $Y=35445
X655 542 360 1 2 BUFFD2BWP7T $T=424880 27840 1 0 $X=424590 $Y=23630
X656 544 375 1 2 BUFFD2BWP7T $T=445600 27840 1 0 $X=445310 $Y=23630
X657 1 2 DCAP16BWP7T $T=147680 43520 0 0 $X=147390 $Y=43285
X658 1 2 DCAP16BWP7T $T=203120 27840 1 0 $X=202830 $Y=23630
X659 1 2 DCAP16BWP7T $T=216000 20000 0 0 $X=215710 $Y=19765
X660 1 2 DCAP16BWP7T $T=233920 20000 0 0 $X=233630 $Y=19765
X661 1 2 DCAP16BWP7T $T=266400 27840 0 0 $X=266110 $Y=27605
X662 1 2 DCAP16BWP7T $T=287120 43520 0 0 $X=286830 $Y=43285
X663 1 2 DCAP16BWP7T $T=311760 35680 0 0 $X=311470 $Y=35445
X664 1 2 DCAP16BWP7T $T=317920 27840 1 0 $X=317630 $Y=23630
X665 1 2 DCAP16BWP7T $T=329120 43520 1 0 $X=328830 $Y=39310
X666 1 2 DCAP16BWP7T $T=345920 43520 0 0 $X=345630 $Y=43285
X667 1 2 DCAP16BWP7T $T=359360 43520 0 0 $X=359070 $Y=43285
X668 1 2 DCAP16BWP7T $T=371120 35680 0 0 $X=370830 $Y=35445
X669 1 2 DCAP16BWP7T $T=371120 43520 0 0 $X=370830 $Y=43285
X670 1 2 DCAP16BWP7T $T=387360 43520 1 0 $X=387070 $Y=39310
X671 1 2 DCAP16BWP7T $T=389600 27840 1 0 $X=389310 $Y=23630
X672 1 2 DCAP16BWP7T $T=399120 27840 0 0 $X=398830 $Y=27605
X673 1 2 DCAP16BWP7T $T=413120 43520 1 0 $X=412830 $Y=39310
X674 1 2 DCAP16BWP7T $T=420960 35680 0 0 $X=420670 $Y=35445
X675 1 2 DCAP16BWP7T $T=428240 27840 1 0 $X=427950 $Y=23630
X676 1 2 DCAP16BWP7T $T=455120 35680 1 0 $X=454830 $Y=31470
X677 1 2 DCAP16BWP7T $T=455120 43520 1 0 $X=454830 $Y=39310
X678 1 2 DCAP16BWP7T $T=464640 20000 0 0 $X=464350 $Y=19765
X679 20 1 2 417 CKND1BWP7T $T=38480 27840 1 0 $X=38190 $Y=23630
X680 418 1 2 85 CKND1BWP7T $T=79920 35680 1 0 $X=79630 $Y=31470
X681 275 1 2 504 CKND1BWP7T $T=265280 35680 1 180 $X=263310 $Y=35445
X682 273 1 2 512 CKND1BWP7T $T=292720 35680 1 180 $X=290750 $Y=35445
X683 301 1 2 302 BUFFD3BWP7T $T=308960 20000 0 0 $X=308670 $Y=19765
X684 518 1 2 315 BUFFD3BWP7T $T=320720 20000 0 0 $X=320430 $Y=19765
X685 519 1 2 316 BUFFD3BWP7T $T=320720 27840 0 0 $X=320430 $Y=27605
X686 523 1 2 333 BUFFD3BWP7T $T=348720 27840 1 0 $X=348430 $Y=23630
X687 283 2 507 237 1 NR2D4BWP7T $T=268640 20000 1 180 $X=261630 $Y=19765
X688 3 5 2 1 INVD2BWP7T $T=21120 43520 0 0 $X=20830 $Y=43285
X689 407 4 2 1 INVD2BWP7T $T=23920 27840 1 180 $X=21390 $Y=27605
X690 141 119 2 1 INVD2BWP7T $T=124160 43520 0 180 $X=121630 $Y=39310
X691 458 113 2 1 INVD2BWP7T $T=130880 27840 0 0 $X=130590 $Y=27605
X692 205 194 2 1 INVD2BWP7T $T=192480 27840 0 180 $X=189950 $Y=23630
X693 285 507 2 1 INVD2BWP7T $T=272000 27840 0 180 $X=269470 $Y=23630
X694 297 292 2 1 INVD2BWP7T $T=301120 27840 0 0 $X=300830 $Y=27605
X695 374 377 2 1 INVD2BWP7T $T=446720 43520 1 0 $X=446430 $Y=39310
X696 376 378 2 1 INVD2BWP7T $T=447280 27840 0 0 $X=446990 $Y=27605
X697 379 381 2 1 INVD2BWP7T $T=458480 27840 0 0 $X=458190 $Y=27605
X698 380 382 2 1 INVD2BWP7T $T=459600 43520 0 0 $X=459310 $Y=43285
X699 384 386 2 1 INVD2BWP7T $T=462400 20000 0 0 $X=462110 $Y=19765
X700 389 390 2 1 INVD2BWP7T $T=465760 35680 1 0 $X=465470 $Y=31470
X701 391 393 2 1 INVD2BWP7T $T=467440 43520 1 0 $X=467150 $Y=39310
X702 392 394 2 1 INVD2BWP7T $T=468560 27840 0 0 $X=468270 $Y=27605
X703 524 531 1 2 338 CKXOR2D1BWP7T $T=361600 35680 1 0 $X=361310 $Y=31470
X704 533 529 1 2 342 CKXOR2D1BWP7T $T=377280 35680 1 0 $X=376990 $Y=31470
X705 2 1 DCAP32BWP7T $T=329120 27840 1 0 $X=328830 $Y=23630
X706 2 1 DCAP32BWP7T $T=350960 27840 0 0 $X=350670 $Y=27605
X707 2 1 DCAP32BWP7T $T=429920 35680 1 0 $X=429630 $Y=31470
X708 2 1 DCAP32BWP7T $T=432720 43520 0 0 $X=432430 $Y=43285
X709 520 308 1 2 309 XNR2D1BWP7T $T=314560 43520 1 0 $X=314270 $Y=39310
X710 314 312 1 2 298 XNR2D1BWP7T $T=324640 43520 1 180 $X=319310 $Y=43285
X711 124 134 2 1 CKND2BWP7T $T=112960 35680 0 0 $X=112670 $Y=35445
X712 170 172 2 1 CKND2BWP7T $T=163920 35680 1 0 $X=163630 $Y=31470
X713 366 368 2 1 CKND2BWP7T $T=435520 20000 0 0 $X=435230 $Y=19765
X714 369 370 2 1 CKND2BWP7T $T=438880 27840 1 0 $X=438590 $Y=23630
X715 387 385 2 1 CKND2BWP7T $T=464080 27840 0 180 $X=461550 $Y=23630
X716 396 397 2 1 CKND2BWP7T $T=470800 27840 1 0 $X=470510 $Y=23630
X717 148 1 2 460 CKND0BWP7T $T=127520 27840 1 0 $X=127230 $Y=23630
X718 482 1 2 197 CKND0BWP7T $T=185760 27840 0 0 $X=185470 $Y=27605
X719 283 1 2 287 CKND0BWP7T $T=274240 35680 0 0 $X=273950 $Y=35445
X720 529 2 530 337 336 524 1 AOI22D2BWP7T $T=359920 27840 1 0 $X=359630 $Y=23630
X721 341 2 529 340 524 534 1 AOI22D2BWP7T $T=384000 20000 1 180 $X=376990 $Y=19765
X722 407 1 2 422 CKBD0BWP7T $T=49680 35680 1 0 $X=49390 $Y=31470
X723 196 1 2 474 CKBD0BWP7T $T=184080 27840 1 180 $X=181550 $Y=27605
X724 6 2 407 8 1 NR2D1BWP7T $T=22240 20000 0 0 $X=21950 $Y=19765
X725 26 2 28 417 1 NR2D1BWP7T $T=40160 27840 1 0 $X=39870 $Y=23630
X726 59 2 427 15 1 NR2D1BWP7T $T=58080 35680 1 180 $X=55550 $Y=35445
X727 67 2 86 440 1 NR2D1BWP7T $T=79920 43520 0 0 $X=79630 $Y=43285
X728 66 2 441 440 1 NR2D1BWP7T $T=84400 35680 1 180 $X=81870 $Y=35445
X729 141 2 150 461 1 NR2D1BWP7T $T=127520 43520 1 0 $X=127230 $Y=39310
X730 165 2 466 156 1 NR2D1BWP7T $T=147680 20000 1 180 $X=145150 $Y=19765
X731 458 2 167 468 1 NR2D1BWP7T $T=147680 27840 0 0 $X=147390 $Y=27605
X732 180 2 182 184 1 NR2D1BWP7T $T=173440 35680 0 0 $X=173150 $Y=35445
X733 197 2 475 202 1 NR2D1BWP7T $T=184640 35680 1 0 $X=184350 $Y=31470
X734 208 2 490 202 1 NR2D1BWP7T $T=196400 20000 0 0 $X=196110 $Y=19765
X735 208 2 480 497 1 NR2D1BWP7T $T=212080 27840 0 0 $X=211790 $Y=27605
X736 263 2 501 256 1 NR2D1BWP7T $T=241200 43520 1 180 $X=238670 $Y=43285
X737 275 2 497 270 1 NR2D1BWP7T $T=260800 27840 1 180 $X=258270 $Y=27605
X738 429 54 57 55 2 1 423 NR4D1BWP7T $T=57520 43520 0 180 $X=51630 $Y=39310
X739 68 70 424 9 2 1 66 NR4D1BWP7T $T=65360 35680 1 180 $X=59470 $Y=35445
X740 439 437 32 430 2 1 435 NR4D1BWP7T $T=70960 27840 1 180 $X=65070 $Y=27605
X741 188 184 476 473 2 1 474 NR4D1BWP7T $T=179040 27840 1 180 $X=173150 $Y=27605
X742 181 180 186 479 2 1 190 NR4D1BWP7T $T=174560 43520 1 0 $X=174270 $Y=39310
X743 195 193 484 481 2 1 204 NR4D1BWP7T $T=182960 35680 0 0 $X=182670 $Y=35445
X744 207 484 202 208 2 1 209 NR4D1BWP7T $T=190800 43520 1 0 $X=190510 $Y=39310
X745 215 202 203 488 2 1 196 NR4D1BWP7T $T=199200 35680 1 180 $X=193310 $Y=35445
X746 212 211 487 491 2 1 216 NR4D1BWP7T $T=193600 43520 0 0 $X=193310 $Y=43285
X747 496 224 494 218 2 1 487 NR4D1BWP7T $T=211520 43520 1 180 $X=205630 $Y=43285
X748 183 484 233 236 2 1 235 NR4D1BWP7T $T=215440 35680 0 0 $X=215150 $Y=35445
X749 238 193 237 499 2 1 223 NR4D1BWP7T $T=217120 27840 0 0 $X=216830 $Y=27605
X750 255 256 259 247 2 1 505 NR4D1BWP7T $T=233360 43520 0 0 $X=233070 $Y=43285
X751 495 508 251 476 2 1 505 NR4D1BWP7T $T=247920 27840 0 0 $X=247630 $Y=27605
X752 22 411 24 413 2 1 418 OR4D1BWP7T $T=37920 35680 0 0 $X=37630 $Y=35445
X753 428 91 73 409 2 1 95 OR4D1BWP7T $T=83840 43520 0 0 $X=83550 $Y=43285
X754 409 437 444 96 1 2 98 OA31D0BWP7T $T=86640 43520 1 0 $X=86350 $Y=39310
X755 294 297 293 296 1 2 514 OA31D0BWP7T $T=301120 43520 1 180 $X=296350 $Y=43285
X756 464 2 159 463 113 1 AOI21D2BWP7T $T=139280 27840 1 180 $X=133950 $Y=27605
X757 284 2 476 511 512 1 AOI21D2BWP7T $T=273680 27840 1 0 $X=273390 $Y=23630
X758 5 1 14 20 2 ND2D1BWP7T $T=28960 43520 0 0 $X=28670 $Y=43285
X759 21 1 23 416 2 ND2D1BWP7T $T=37920 43520 1 0 $X=37630 $Y=39310
X760 21 1 415 25 2 ND2D1BWP7T $T=37920 43520 0 0 $X=37630 $Y=43285
X761 30 1 414 20 2 ND2D1BWP7T $T=41840 35680 0 180 $X=39310 $Y=31470
X762 33 1 35 19 2 ND2D1BWP7T $T=42400 35680 0 0 $X=42110 $Y=35445
X763 25 1 36 20 2 ND2D1BWP7T $T=42960 43520 0 0 $X=42670 $Y=43285
X764 23 1 40 414 2 ND2D1BWP7T $T=47440 43520 0 180 $X=44910 $Y=39310
X765 27 1 43 416 2 ND2D1BWP7T $T=45760 43520 0 0 $X=45470 $Y=43285
X766 16 1 45 33 2 ND2D1BWP7T $T=47440 35680 1 0 $X=47150 $Y=31470
X767 19 1 48 416 2 ND2D1BWP7T $T=47440 43520 1 0 $X=47150 $Y=39310
X768 27 1 50 51 2 ND2D1BWP7T $T=49120 43520 0 0 $X=48830 $Y=43285
X769 33 1 52 422 2 ND2D1BWP7T $T=50240 27840 0 0 $X=49950 $Y=27605
X770 422 1 53 51 2 ND2D1BWP7T $T=53600 43520 1 180 $X=51070 $Y=43285
X771 36 1 424 23 2 ND2D1BWP7T $T=51920 35680 0 0 $X=51630 $Y=35445
X772 47 1 63 422 2 ND2D1BWP7T $T=58080 27840 0 0 $X=57790 $Y=27605
X773 63 1 435 23 2 ND2D1BWP7T $T=70400 35680 0 180 $X=67870 $Y=31470
X774 84 1 70 427 2 ND2D1BWP7T $T=80480 43520 1 0 $X=80190 $Y=39310
X775 107 1 448 104 2 ND2D1BWP7T $T=96160 43520 1 180 $X=93630 $Y=43285
X776 108 1 111 113 2 ND2D1BWP7T $T=98400 43520 0 0 $X=98110 $Y=43285
X777 112 1 116 452 2 ND2D1BWP7T $T=100640 43520 0 0 $X=100350 $Y=43285
X778 124 1 127 452 2 ND2D1BWP7T $T=106800 43520 0 0 $X=106510 $Y=43285
X779 148 1 142 139 2 ND2D1BWP7T $T=126400 35680 1 180 $X=123870 $Y=35445
X780 119 1 149 148 2 ND2D1BWP7T $T=124720 43520 1 0 $X=124430 $Y=39310
X781 143 1 144 452 2 ND2D1BWP7T $T=124720 43520 0 0 $X=124430 $Y=43285
X782 143 1 107 139 2 ND2D1BWP7T $T=134800 43520 1 180 $X=132270 $Y=43285
X783 467 1 110 454 2 ND2D1BWP7T $T=145440 35680 0 180 $X=142910 $Y=31470
X784 465 1 468 165 2 ND2D1BWP7T $T=147680 20000 0 0 $X=147390 $Y=19765
X785 169 1 128 170 2 ND2D1BWP7T $T=149360 43520 1 0 $X=149070 $Y=39310
X786 467 1 171 156 2 ND2D1BWP7T $T=151040 20000 0 0 $X=150750 $Y=19765
X787 172 1 145 169 2 ND2D1BWP7T $T=153840 43520 0 180 $X=151310 $Y=39310
X788 482 1 486 206 2 ND2D1BWP7T $T=190800 27840 0 0 $X=190510 $Y=27605
X789 495 1 225 480 2 ND2D1BWP7T $T=213200 35680 0 180 $X=210670 $Y=31470
X790 242 1 227 241 2 ND2D1BWP7T $T=224960 35680 1 180 $X=222430 $Y=35445
X791 503 1 483 243 2 ND2D1BWP7T $T=230560 27840 1 180 $X=228030 $Y=27605
X792 250 1 243 239 2 ND2D1BWP7T $T=230560 35680 1 180 $X=228030 $Y=35445
X793 242 1 248 252 2 ND2D1BWP7T $T=228880 35680 1 0 $X=228590 $Y=31470
X794 504 1 232 253 2 ND2D1BWP7T $T=235040 43520 0 180 $X=232510 $Y=39310
X795 254 1 502 258 2 ND2D1BWP7T $T=237280 43520 0 180 $X=234750 $Y=39310
X796 250 1 260 262 2 ND2D1BWP7T $T=241200 43520 0 180 $X=238670 $Y=39310
X797 250 1 509 268 2 ND2D1BWP7T $T=250720 35680 0 0 $X=250430 $Y=35445
X798 273 1 503 268 2 ND2D1BWP7T $T=261360 35680 1 180 $X=258830 $Y=35445
X799 294 1 515 516 2 ND2D1BWP7T $T=306160 43520 1 0 $X=305870 $Y=39310
X800 14 1 12 410 2 411 11 OAI211D1BWP7T $T=29520 35680 1 180 $X=25870 $Y=35445
X801 450 2 446 94 89 1 106 NR4D2BWP7T $T=96160 20000 1 180 $X=82990 $Y=19765
X802 505 2 194 236 223 1 228 NR4D2BWP7T $T=238960 27840 0 180 $X=225790 $Y=23630
X803 511 2 279 272 1 NR2XD0BWP7T $T=271440 35680 0 180 $X=268910 $Y=31470
X804 37 1 31 415 414 29 2 ND4D1BWP7T $T=45200 43520 0 180 $X=40990 $Y=39310
X805 35 1 414 41 12 420 2 ND4D1BWP7T $T=44640 35680 0 0 $X=44350 $Y=35445
X806 50 1 65 436 429 82 2 ND4D1BWP7T $T=68720 43520 0 0 $X=68430 $Y=43285
X807 79 1 441 429 85 443 2 ND4D1BWP7T $T=83280 35680 1 0 $X=82990 $Y=31470
X808 226 1 496 219 228 230 2 ND4D1BWP7T $T=211520 43520 1 0 $X=211230 $Y=39310
X809 226 1 234 500 501 190 2 ND4D1BWP7T $T=217120 43520 0 0 $X=216830 $Y=43285
X810 465 156 455 128 121 1 2 OAI31D1BWP7T $T=136480 27840 0 180 $X=132270 $Y=23630
X811 292 291 513 511 290 1 2 OAI31D1BWP7T $T=281520 27840 1 180 $X=277310 $Y=27605
X812 424 1 2 423 46 412 38 NR4D0BWP7T $T=54720 27840 1 0 $X=54430 $Y=23630
X813 62 1 2 423 15 425 28 NR4D0BWP7T $T=58080 27840 1 180 $X=54430 $Y=27605
X814 78 1 2 409 24 438 433 NR4D0BWP7T $T=70400 35680 1 180 $X=66750 $Y=35445
X815 203 1 2 198 197 200 184 NR4D0BWP7T $T=186320 43520 1 180 $X=182670 $Y=43285
X816 493 1 2 231 499 489 193 NR4D0BWP7T $T=214320 27840 1 0 $X=214030 $Y=23630
X817 502 1 2 240 236 500 233 NR4D0BWP7T $T=222720 43520 0 180 $X=219070 $Y=39310
X818 249 1 2 203 247 245 494 NR4D0BWP7T $T=229440 43520 1 180 $X=225790 $Y=43285
X819 61 26 2 431 1 NR2D2BWP7T $T=59200 20000 0 0 $X=58910 $Y=19765
X820 101 453 2 99 1 NR2D2BWP7T $T=96720 27840 0 0 $X=96430 $Y=27605
X821 270 293 2 240 1 NR2D2BWP7T $T=294960 43520 0 180 $X=290750 $Y=39310
X822 297 516 2 506 1 NR2D2BWP7T $T=307840 27840 0 180 $X=303630 $Y=23630
X823 438 43 81 79 2 1 76 AN4D1BWP7T $T=73200 43520 0 180 $X=68990 $Y=39310
X824 425 1 2 426 BUFFD0BWP7T $T=52480 27840 0 0 $X=52190 $Y=27605
X825 439 1 2 83 BUFFD0BWP7T $T=70960 27840 0 0 $X=70670 $Y=27605
X826 12 1 48 53 58 428 2 ND4D0BWP7T $T=53600 43520 0 0 $X=53310 $Y=43285
X827 65 1 63 23 45 432 2 ND4D0BWP7T $T=63680 35680 0 180 $X=60030 $Y=31470
X828 52 1 90 85 427 88 2 ND4D0BWP7T $T=86640 43520 0 180 $X=82990 $Y=39310
X829 84 1 442 93 441 444 2 ND4D0BWP7T $T=84400 35680 0 0 $X=84110 $Y=35445
X830 192 1 214 489 490 491 2 ND4D0BWP7T $T=195280 27840 1 0 $X=194990 $Y=23630
X831 221 1 219 220 213 472 2 ND4D0BWP7T $T=209280 35680 1 180 $X=205630 $Y=35445
X832 449 445 447 2 1 NR2D1P5BWP7T $T=94480 35680 0 180 $X=90270 $Y=31470
X833 449 459 101 2 1 NR2D1P5BWP7T $T=123600 27840 1 0 $X=123310 $Y=23630
X834 178 169 177 2 1 NR2D1P5BWP7T $T=167840 43520 1 0 $X=167550 $Y=39310
X835 484 201 485 2 1 NR2D1P5BWP7T $T=189120 43520 0 180 $X=184910 $Y=39310
X836 279 508 507 2 1 NR2D1P5BWP7T $T=265840 27840 1 0 $X=265550 $Y=23630
X837 294 299 298 2 1 NR2D1P5BWP7T $T=300560 43520 1 0 $X=300270 $Y=39310
X838 287 506 504 2 1 488 OA21D0BWP7T $T=268640 35680 1 180 $X=264990 $Y=35445
X839 483 1 482 192 2 473 IND3D0BWP7T $T=184080 27840 0 180 $X=180430 $Y=23630
X840 483 1 482 192 2 199 IND3D0BWP7T $T=188560 27840 0 180 $X=184910 $Y=23630
X841 433 1 406 69 72 2 NR3D1BWP7T $T=62560 43520 1 0 $X=62270 $Y=39310
X842 459 1 136 135 147 2 NR3D1BWP7T $T=130320 35680 0 180 $X=125550 $Y=31470
X843 493 1 483 486 222 2 NR3D1BWP7T $T=205920 27840 0 0 $X=205630 $Y=27605
X844 208 1 483 498 229 2 NR3D1BWP7T $T=216000 20000 1 180 $X=211230 $Y=19765
X845 180 1 475 477 481 189 2 IND4D0BWP7T $T=175680 35680 0 0 $X=175390 $Y=35445
X846 126 1 133 131 450 104 2 IND4D1BWP7T $T=113520 43520 1 180 $X=108750 $Y=43285
X847 497 1 248 246 485 244 2 IND4D1BWP7T $T=230000 43520 0 180 $X=225230 $Y=39310
X848 231 1 248 258 498 254 2 IND4D1BWP7T $T=237840 27840 1 180 $X=233070 $Y=27605
X849 29 432 431 34 2 1 434 OR4D0BWP7T $T=63680 35680 1 0 $X=63390 $Y=31470
X850 176 177 137 2 1 INR2D2BWP7T $T=165040 43520 0 0 $X=164750 $Y=43285
X851 289 282 290 2 1 INR2D2BWP7T $T=277600 43520 1 0 $X=277310 $Y=39310
X852 4 2 406 1 3 NR2XD1BWP7T $T=21120 35680 1 0 $X=20830 $Y=31470
X853 3 2 409 1 410 NR2XD1BWP7T $T=24480 27840 0 0 $X=24190 $Y=27605
X854 13 2 15 1 410 NR2XD1BWP7T $T=27280 20000 0 0 $X=26990 $Y=19765
X855 17 2 16 1 8 NR2XD1BWP7T $T=31200 35680 0 180 $X=26990 $Y=31470
X856 417 2 38 1 39 NR2XD1BWP7T $T=42960 20000 0 0 $X=42670 $Y=19765
X857 26 2 46 1 410 NR2XD1BWP7T $T=46880 20000 0 0 $X=46590 $Y=19765
X858 419 2 56 1 39 NR2XD1BWP7T $T=50800 20000 0 0 $X=50510 $Y=19765
X859 421 2 54 1 410 NR2XD1BWP7T $T=54720 27840 0 180 $X=50510 $Y=23630
X860 61 2 60 1 39 NR2XD1BWP7T $T=59200 20000 1 180 $X=54990 $Y=19765
X861 431 2 80 1 60 NR2XD1BWP7T $T=73200 20000 1 180 $X=68990 $Y=19765
X862 447 2 102 1 451 NR2XD1BWP7T $T=91680 35680 0 0 $X=91390 $Y=35445
X863 110 2 114 1 451 NR2XD1BWP7T $T=98960 35680 0 0 $X=98670 $Y=35445
X864 456 2 115 1 453 NR2XD1BWP7T $T=103440 27840 0 180 $X=99230 $Y=23630
X865 449 2 118 1 456 NR2XD1BWP7T $T=105680 20000 1 180 $X=101470 $Y=19765
X866 128 2 123 1 110 NR2XD1BWP7T $T=109040 35680 0 180 $X=104830 $Y=31470
X867 126 2 457 1 445 NR2XD1BWP7T $T=109040 35680 1 180 $X=104830 $Y=35445
X868 101 2 125 1 451 NR2XD1BWP7T $T=106240 27840 0 0 $X=105950 $Y=27605
X869 456 2 126 1 451 NR2XD1BWP7T $T=107360 20000 0 0 $X=107070 $Y=19765
X870 128 2 129 1 132 NR2XD1BWP7T $T=109040 27840 1 0 $X=108750 $Y=23630
X871 451 2 130 1 134 NR2XD1BWP7T $T=109040 35680 0 0 $X=108750 $Y=35445
X872 449 2 135 1 132 NR2XD1BWP7T $T=111280 20000 0 0 $X=110990 $Y=19765
X873 458 2 136 1 132 NR2XD1BWP7T $T=115200 27840 1 180 $X=110990 $Y=27605
X874 145 2 140 1 132 NR2XD1BWP7T $T=125840 35680 0 180 $X=121630 $Y=31470
X875 460 2 138 1 458 NR2XD1BWP7T $T=126960 27840 1 180 $X=122750 $Y=27605
X876 460 2 146 1 449 NR2XD1BWP7T $T=128080 20000 1 180 $X=123870 $Y=19765
X877 152 2 151 1 136 NR2XD1BWP7T $T=130880 43520 1 180 $X=126670 $Y=43285
X878 460 2 155 1 453 NR2XD1BWP7T $T=131440 35680 1 0 $X=131150 $Y=31470
X879 468 2 148 1 156 NR2XD1BWP7T $T=143200 27840 0 180 $X=138990 $Y=23630
X880 469 2 176 1 170 NR2XD1BWP7T $T=170080 35680 1 180 $X=165870 $Y=35445
X881 270 2 235 1 507 NR2XD1BWP7T $T=256880 27840 0 180 $X=252670 $Y=23630
X882 275 2 223 1 279 NR2XD1BWP7T $T=259680 27840 1 0 $X=259390 $Y=23630
X883 275 2 180 1 284 NR2XD1BWP7T $T=271440 43520 0 180 $X=267230 $Y=39310
X884 271 2 233 1 511 NR2XD1BWP7T $T=276480 20000 1 180 $X=272270 $Y=19765
X885 512 2 203 1 280 NR2XD1BWP7T $T=279840 35680 1 180 $X=275630 $Y=35445
X886 515 2 239 1 297 NR2XD1BWP7T $T=302800 35680 1 180 $X=298590 $Y=35445
X887 516 2 510 1 292 NR2XD1BWP7T $T=312320 27840 1 180 $X=308110 $Y=27605
X888 80 2 406 437 97 443 1 INR4D2BWP7T $T=79920 27840 1 0 $X=79630 $Y=23630
X889 206 2 194 478 185 471 1 INR4D2BWP7T $T=188560 20000 1 180 $X=173710 $Y=19765
X890 14 1 12 11 10 410 2 OAI211D2BWP7T $T=30640 43520 0 180 $X=24190 $Y=39310
X891 31 1 414 39 42 17 2 OAI211D2BWP7T $T=40720 27840 0 0 $X=40430 $Y=27605
X892 120 1 151 461 158 453 2 OAI211D2BWP7T $T=130880 43520 1 0 $X=130590 $Y=39310
X893 241 1 239 482 2 CKND2D0BWP7T $T=222160 35680 0 180 $X=219630 $Y=31470
X894 454 452 459 153 1 2 462 AO211D0BWP7T $T=128640 35680 0 0 $X=128350 $Y=35445
X895 261 510 497 272 1 2 492 AO211D0BWP7T $T=258560 35680 0 180 $X=254350 $Y=31470
X896 448 2 445 109 454 452 1 AOI211D2BWP7T $T=93920 43520 1 0 $X=93630 $Y=39310
X897 257 2 187 221 506 261 1 AOI211D2BWP7T $T=233360 35680 1 0 $X=233070 $Y=31470
X898 265 2 256 267 510 504 1 AOI211D2BWP7T $T=250160 43520 1 0 $X=249870 $Y=39310
X899 13 2 32 417 1 NR2D3BWP7T $T=37920 20000 0 0 $X=37630 $Y=19765
X900 447 2 117 453 1 NR2D3BWP7T $T=99520 35680 1 0 $X=99230 $Y=31470
X901 141 2 160 134 1 NR2D3BWP7T $T=134800 43520 0 0 $X=134510 $Y=43285
X902 132 2 168 453 1 NR2D3BWP7T $T=153280 35680 0 180 $X=147950 $Y=31470
X903 283 2 288 511 1 NR2D3BWP7T $T=276480 35680 0 180 $X=271150 $Y=31470
X904 512 2 184 279 1 NR2D3BWP7T $T=277040 43520 0 180 $X=271710 $Y=39310
X905 275 2 282 271 1 NR2D3BWP7T $T=298320 20000 1 180 $X=292990 $Y=19765
X906 515 2 268 292 1 NR2D3BWP7T $T=308400 35680 0 180 $X=303070 $Y=31470
X907 517 2 273 300 1 NR2D3BWP7T $T=314000 43520 0 180 $X=308670 $Y=39310
X908 27 25 1 2 34 AN2D1BWP7T $T=40160 43520 0 0 $X=39870 $Y=43285
X909 416 422 1 2 59 AN2D1BWP7T $T=51920 35680 1 0 $X=51630 $Y=31470
X910 422 25 1 2 62 AN2D1BWP7T $T=64800 27840 1 180 $X=61710 $Y=27605
X911 165 467 1 2 175 AN2D1BWP7T $T=167280 20000 1 180 $X=164190 $Y=19765
X912 170 174 1 2 139 AN2D1BWP7T $T=167840 43520 0 180 $X=164750 $Y=39310
X913 8 410 408 1 2 ND2D2BWP7T $T=29520 27840 0 180 $X=25310 $Y=23630
X914 122 121 119 1 2 ND2D2BWP7T $T=107920 43520 0 180 $X=103710 $Y=39310
X915 174 453 172 1 2 ND2D2BWP7T $T=156080 35680 1 180 $X=151870 $Y=35445
X916 173 132 175 1 2 ND2D2BWP7T $T=164480 27840 1 0 $X=164190 $Y=23630
X917 506 279 291 1 2 ND2D2BWP7T $T=282080 35680 0 180 $X=277870 $Y=31470
X918 294 270 506 1 2 ND2D2BWP7T $T=292160 27840 1 0 $X=291870 $Y=23630
X919 294 283 510 1 2 ND2D2BWP7T $T=301120 27840 1 180 $X=296910 $Y=27605
X920 281 275 300 1 2 ND2D2BWP7T $T=308960 43520 1 180 $X=304750 $Y=43285
X921 466 139 1 117 161 2 AOI21D1BWP7T $T=141520 43520 0 180 $X=137870 $Y=39310
X922 53 64 50 37 430 1 2 ND4D2BWP7T $T=56960 43520 0 0 $X=56670 $Y=43285
X923 266 269 509 503 218 1 2 ND4D2BWP7T $T=251280 43520 0 0 $X=250990 $Y=43285
X924 71 2 73 422 1 436 25 AOI211D1BWP7T $T=64240 43520 0 0 $X=63950 $Y=43285
X925 227 2 213 223 1 INR2D1BWP7T $T=212640 35680 1 180 $X=209550 $Y=35445
X926 99 94 2 1 CKBD2BWP7T $T=91680 27840 1 180 $X=88030 $Y=27605
X928 319 327 323 332 2 1 545 DFCND1BWP7T $T=339200 43520 1 0 $X=338910 $Y=39310
X929 319 539 323 336 2 1 530 DFCND1BWP7T $T=399120 27840 1 180 $X=385950 $Y=27605
X930 319 541 323 341 2 1 534 DFCND1BWP7T $T=404720 20000 1 180 $X=391550 $Y=19765
X931 528 522 467 1 2 XNR2D2BWP7T $T=362160 20000 1 180 $X=355150 $Y=19765
X932 319 358 323 362 546 1 2 DFCND2BWP7T $T=418160 43520 0 0 $X=417870 $Y=43285
X933 319 328 323 318 2 1 520 DFCND0BWP7T $T=345920 43520 1 180 $X=332750 $Y=43285
X934 319 535 323 532 2 1 531 DFCND0BWP7T $T=387360 43520 0 180 $X=374190 $Y=39310
X935 319 537 323 527 2 1 547 DFCND0BWP7T $T=389600 27840 0 180 $X=376430 $Y=23630
X936 319 536 323 538 2 1 533 DFCND0BWP7T $T=380080 35680 0 0 $X=379790 $Y=35445
X937 353 347 345 336 343 341 2 540 1 OA222D0BWP7T $T=405840 43520 1 180 $X=399390 $Y=43285
X938 208 2 282 1 277 281 262 AOI211XD1BWP7T $T=268640 43520 1 180 $X=261630 $Y=43285
X939 305 307 1 2 INVD2P5BWP7T $T=315120 27840 1 0 $X=314830 $Y=23630
X940 317 321 1 2 INVD2P5BWP7T $T=334160 20000 0 0 $X=333870 $Y=19765
X941 324 326 1 2 INVD2P5BWP7T $T=339200 20000 0 0 $X=338910 $Y=19765
X942 329 330 1 2 INVD2P5BWP7T $T=346480 20000 0 0 $X=346190 $Y=19765
X943 372 373 1 2 INVD2P5BWP7T $T=442800 20000 0 0 $X=442510 $Y=19765
X944 383 388 1 2 INVD2P5BWP7T $T=461840 35680 0 0 $X=461550 $Y=35445
X945 395 398 1 2 INVD2P5BWP7T $T=470240 43520 1 0 $X=469950 $Y=39310
X946 347 348 1 345 532 343 344 2 535 OAI222D2BWP7T $T=391840 43520 1 180 $X=381470 $Y=43285
X947 347 350 1 345 538 343 532 2 536 OAI222D2BWP7T $T=403040 35680 1 180 $X=392670 $Y=35445
X948 347 354 1 345 335 343 538 2 537 OAI222D2BWP7T $T=407520 43520 0 180 $X=397150 $Y=39310
X949 461 2 1 467 108 NR2D2P5BWP7T $T=139840 27840 0 0 $X=139550 $Y=27605
X950 165 2 1 173 454 NR2D2P5BWP7T $T=151600 27840 1 0 $X=151310 $Y=23630
X951 275 2 1 280 231 NR2D2P5BWP7T $T=261360 27840 0 0 $X=261070 $Y=27605
X952 283 2 1 293 295 NR2D2P5BWP7T $T=299440 35680 0 180 $X=294110 $Y=31470
X953 273 239 1 2 265 CKAN2D1BWP7T $T=259120 35680 1 180 $X=256030 $Y=35445
X954 420 2 424 34 77 1 NR3D2BWP7T $T=60320 27840 1 0 $X=60030 $Y=23630
X955 164 141 459 163 2 1 IAO21D2BWP7T $T=146000 43520 1 180 $X=140670 $Y=43285
X956 465 101 454 1 2 ND2D1P5BWP7T $T=147680 27840 1 0 $X=147390 $Y=23630
X957 510 284 291 1 2 ND2D1P5BWP7T $T=278720 27840 1 0 $X=278430 $Y=23630
X958 202 213 214 210 1 2 486 IIND4D1BWP7T $T=193040 27840 0 0 $X=192750 $Y=27605
X959 239 271 1 2 INVD1P5BWP7T $T=289920 35680 1 0 $X=289630 $Y=31470
X960 155 2 146 454 1 162 157 AOI211XD2BWP7T $T=147680 35680 1 180 $X=134510 $Y=35445
X961 461 2 1 122 465 NR2XD2BWP7T $T=133120 20000 0 0 $X=132830 $Y=19765
X962 173 2 1 124 468 NR2XD2BWP7T $T=156640 27840 1 180 $X=149630 $Y=27605
X963 271 2 1 193 507 NR2XD2BWP7T $T=255200 20000 1 180 $X=248190 $Y=19765
X964 250 242 202 1 2 AN2D2BWP7T $T=233920 20000 1 180 $X=229710 $Y=19765
X965 406 7 9 1 2 IND2D2BWP7T $T=26160 35680 1 180 $X=21390 $Y=35445
X966 275 2 283 1 263 NR2XD3BWP7T $T=280960 43520 1 180 $X=272270 $Y=43285
X967 454 1 467 2 463 OR2D0BWP7T $T=146000 27840 0 180 $X=142910 $Y=23630
X968 367 364 322 1 2 INR2XD4BWP7T $T=440000 27840 1 180 $X=426830 $Y=27605
X969 367 365 314 1 2 INR2XD4BWP7T $T=440560 43520 0 180 $X=427390 $Y=39310
X970 367 371 333 1 2 INR2XD4BWP7T $T=447280 35680 1 180 $X=434110 $Y=35445
X971 421 1 419 2 44 OR2D1BWP7T $T=50240 27840 0 180 $X=47150 $Y=23630
.ENDS
***************************************
.SUBCKT clefia_128 VDD VSS clk p<69> p<72> p<67> k<110> reset_n p<27> p<24> p<22> p<28> p<53> p<25> k<124> k<60> p<57> k<28> p<59> k<104>
+ p<33> p<26> p<46> p<39> k<102> k<88> p<4> k<103> k<94> done k<100> p<2> p<19> k<101> k<66> k<58> k<45> k<41> k<59> k<46>
+ k<52> k<36> k<25> k<33> k<21> k<23> k<7> k<27> k<14> k<35> k<24> k<9> k<1> k<2> c<93> k<12> c<124> k<0> k<11> c<127>
+ c<121> k<6> k<4> c<125> c<77> c<30> c<36> c<37> c<32> c<33> c<31> c<29> k<111> p<70> p<71> p<73> p<74> p<75> p<76> p<77>
+ p<78> p<79> p<80> p<81> p<82> p<83> p<84> p<85> p<86> p<87> p<88> p<89> p<90> p<91> p<92> p<93> p<94> p<95> p<96> p<97>
+ p<98> p<99> p<100> p<101> p<102> p<103> p<104> p<105> p<106> p<107> p<108> p<109> p<110> p<111> p<112> p<113> p<114> p<115> p<116> p<117>
+ p<118> p<119> p<120> p<121> p<122> p<123> p<124> p<125> p<126> p<127> start p<29> p<30> p<31> p<32> p<34> p<35> p<36> p<37> p<38>
+ p<40> p<41> p<42> p<43> p<44> p<45> p<47> p<48> p<49> p<50> p<51> p<52> p<54> p<55> p<56> p<58> p<60> p<61> p<62> p<63>
+ p<64> p<65> p<66> p<68> k<105> k<106> k<107> k<108> k<109> k<112> k<113> k<114> k<115> k<116> k<117> k<118> k<119> k<120> k<121> k<122>
+ k<123> k<125> k<126> k<127> p<0> p<1> p<3> p<5> p<6> p<7> p<8> p<9> p<10> p<11> p<12> p<13> p<14> p<15> p<16> p<17>
+ p<18> p<20> p<21> p<23> k<51> k<53> k<54> k<55> k<56> k<57> k<61> k<62> k<63> k<64> k<65> k<67> k<68> k<69> k<70> k<71>
+ k<72> k<73> k<74> k<75> k<76> k<77> k<78> k<79> k<80> k<81> k<82> k<83> k<84> k<85> k<86> k<87> k<89> k<90> k<91> k<92>
+ k<93> k<95> k<96> k<97> k<98> k<99> c<14> k<29> k<30> k<31> k<32> k<34> k<37> k<38> k<39> k<40> k<42> k<43> k<44> k<47>
+ k<48> k<49> k<50> k<3> k<5> k<8> k<10> k<13> k<15> k<16> k<17> k<18> k<19> k<20> k<22> k<26> c<82> c<83> c<84> c<85>
+ c<86> c<87> c<88> c<89> c<90> c<91> c<92> c<94> c<95> c<96> c<97> c<98> c<99> c<100> c<101> c<102> c<103> c<104> c<105> c<106>
+ c<107> c<108> c<109> c<110> c<111> c<112> c<113> c<114> c<115> c<116> c<117> c<118> c<119> c<120> c<122> c<123> c<126> c<35> c<38> c<39>
+ c<40> c<41> c<42> c<43> c<44> c<45> c<46> c<47> c<48> c<49> c<50> c<51> c<52> c<53> c<54> c<55> c<56> c<57> c<58> c<59>
+ c<60> c<61> c<62> c<63> c<64> c<65> c<66> c<67> c<68> c<69> c<70> c<71> c<72> c<73> c<74> c<75> c<76> c<78> c<79> c<80>
+ c<81> c<0> c<1> c<2> c<3> c<4> c<5> c<6> c<7> c<8> c<9> c<10> c<11> c<12> c<13> c<15> c<16> c<17> c<18> c<19>
+ c<20> c<21> c<22> c<23> c<24> c<25> c<26> c<27> c<28> c<34>
** N=2740 EP=390 IP=6596 FDC=74353
X0 VSS VDD 52 4 clk 7 54 5 6 14 1874 10 1862 1860 8 9 1861 1865 25 13
+ 12 17 11 28 1863 1871 15 1864 1887 16 1495 18 1866 19 1867 21 23 30 20 22
+ 1869 1868 24 1870 40 27 26 29 31 34 35 1872 39 33 1875 1876 36 1873 37 1879
+ 1878 38 1877 41 42 43 1881 1886 1880 1885 32 1882 44 1883 1884 1496 45 46 1889 164
+ 47 1888 48 49 51 53 1890 50 115 55 58 109 1891 56 1899 57 1941 97 1944 1966
+ 59 1892 1896 60 1894 61 1898 1897 1895 1903 1956 62 1906 1905 1910 63 1904 1923 64 1900
+ 1940 1909 1908 1901 67 81 65 1917 1907 74 68 66 1919 1497 93 69 1928 1925 70 1902
+ 1926 71 79 72 1912 1911 73 1953 75 1922 1915 1914 1918 1916 1936 1947 1924 78 1920 76
+ 77 1921 1893 1929 1963 85 1932 1939 1930 92 1931 1927 84 1933 83 82 1938 90 1935 1934
+ 80 1913 87 88 1937 86 1960 1948 1945 89 1946 1943 91 1949 94 1954 100 95 96 1952
+ 107 1951 1950 1957 1958 103 1942 98 99 101 1959 1955 105 106 104 1961 1964 1962 111 108
+ 465 start 1970 110 1967 113 1969 1968 119 114 120 1965 116 1973 1974 1972 117 1971 1976 1985
+ 1975 121 1977 127 118 122 561 1978 193 915 146 1980 124 125 126 1988 1982 129 131 1984
+ 128 311 2002 130 168 185 2005 132 1987 p<80> 136 133 p<112> 1986 349 135 p<104> 1979 p<76> 123
+ 137 138 360 p<108> 1995 134 932 139 2011 p<115> 1992 1989 1990 1498 140 1991 141 147 142 919
+ 143 112 144 145 p<83> 1983 1993 2018 p<69> 2009 p<122> 1994 p<90> 154 152 1996 1997 149 1647 376
+ 150 153 151 p<111> 1999 p<125> 1998 155 156 2001 569 157 2000 160 p<93> 183 927 159 928 163
+ 737 162 p<67> 165 166 p<99> 2006 331 p<127> p<113> 2003 2007 p<81> 548 169 314 170 p<86> 174 171
+ p<120> p<88> p<118> 2008 2004 939 p<75> 176 573 173 p<78> 175 p<79> 2013 p<107> 172 2015 161 p<95> 2010
+ c<93> 354 178 179 181 p<102> 180 k<110> 578 182 2012 357 reset_n p<110> 2014 184 364 282 2016 p<70>
+ p<96> 186 187 188 p<82> p<71> p<85> 2017 p<92> 593 190 192 189 371 p<114> 191 194 k<127> p<77> 2019
+ p<117> done p<106> p<103> 195 p<124> p<123> p<109> 592 197 196 p<87> 1294 p<121> p<91> 1981 p<74> 2021 p<119> p<84>
+ p<89> p<94> p<97> 588 2020 p<126> k<125> k<111> p<105> c<92> p<101> p<98> p<73> p<100> p<72> p<116>
+ ICV_16 $T=0 0 0 0 $X=2540 $Y=415600
X1 VSS VDD 4 200 199 12 5 202 203 6 2022 10 1860 212 8 2028 228 2035 2090 2088
+ 253 2027 2030 204 2024 11 201 222 1865 1862 205 2025 1890 1495 1861 206 208 213 207 13
+ 210 2058 209 226 9 28 2026 1863 2023 2029 2034 15 14 2051 1888 255 2036 2033 2031 16
+ 240 2038 1562 2068 1866 211 2032 244 2044 19 46 216 2043 214 20 215 18 1869 2037 1558
+ 224 21 22 1496 55 2042 2039 23 1868 1867 220 1559 32 2047 7 25 245 218 2041 2049
+ 219 2048 2045 261 24 1870 2050 1872 26 221 27 2052 40 1873 2054 1883 225 2053 234 252
+ 223 2046 29 2055 1875 2056 2057 242 2060 266 2040 229 33 34 1561 217 230 231 1876 1878
+ 1874 267 31 2079 30 233 2066 35 2061 47 235 2059 2078 37 36 232 1889 38 236 237
+ 241 1879 238 1877 2062 239 227 2063 2074 2064 243 39 2073 41 1880 42 250 43 1881 1882
+ 246 1563 1884 2065 50 247 248 1885 1886 2067 2069 2071 44 249 45 2070 2085 251 2084 2075
+ 2072 48 1887 254 2076 51 49 257 256 2077 263 260 2080 2081 258 2082 53 2086 52 259
+ 2083 262 1564 54 269 264 2087 56 61 265 1892 58 60 2093 1893 268 64 1959 1895 1900
+ 270 62 79 1901 91 271 1902 1897 1955 63 1891 1896 1915 76 67 1916 1899 1907 272 95
+ 68 66 59 1903 2095 1898 1905 1906 1904 70 1911 2089 65 57 1909 69 1913 1910 1497 71
+ 2094 1912 72 75 1965 1918 73 1894 1908 1917 1933 1949 1919 74 1914 1920 82 273 1931 1928
+ 1971 1923 1924 1922 98 1929 78 1926 1921 1925 77 80 1927 1930 81 83 88 102 86 94
+ 274 1938 101 84 1932 1939 93 85 1945 1934 1935 1936 87 275 1943 1942 1940 1937 276 1944
+ 89 97 90 92 1947 1941 1948 96 1950 1946 1952 105 1951 100 2096 1954 99 107 1956 1958
+ 103 1960 2126 104 1957 1953 106 280 2114 2107 1963 1566 2105 281 1966 1976 108 109 149 289
+ 113 1967 2099 110 1968 2120 114 282 284 1974 291 285 2104 2109 115 112 1980 111 116 287
+ 303 2116 2103 128 288 2102 290 283 299 2122 1074 2130 278 193 1979 2108 117 p<65> 119 120
+ 286 2100 2110 2113 292 2111 118 121 2101 123 295 2112 550 296 293 1498 297 194 521 298
+ 2118 2117 300 2119 302 294 1983 301 127 2115 304 129 308 306 305 546 p<30> p<73> 131 2123
+ 307 2124 130 136 2127 185 132 134 309 p<105> 310 135 p<104> 2106 p<98> 2125 126 2128 p<66> p<100>
+ 311 133 137 125 279 2121 528 p<101> 313 172 p<47> 1989 141 139 2097 143 1990 157 145 1998
+ 2129 316 531 142 335 p<68> 1997 314 315 p<29> 2145 2133 312 376 151 146 163 321 162 1647
+ 317 195 942 150 2137 153 154 324 159 152 320 183 2092 322 155 928 323 169 365 p<72>
+ 2143 344 160 382 2136 161 325 p<41> 2135 k<118> 327 164 277 165 330 329 333 168 328 p<56>
+ 2142 2091 331 2144 332 2004 326 564 2140 170 k<86> 2010 p<63> p<22> 762 336 338 181 343 196
+ 340 341 337 176 342 c<79> 345 346 593 2146 339 k<110> 347 350 348 2151 356 362 351 174
+ k<60> 189 180 352 2149 184 355 353 2098 358 489 k<124> p<42> 359 k<99> 361 2148 173 363 2147
+ p<54> 369 2139 2016 589 p<64> 187 p<28> p<52> p<58> 191 188 k<92> 937 2156 2152 p<49> 2131 2134 171
+ 122 p<55> 2157 p<51> 374 k<28> k<47> k<104> 182 2155 k<105> 2138 378 2153 p<61> 379 2141 p<48> 2154 527
+ 2132 p<62> p<40> c<86> p<36> 381 574 384 p<60> 537 p<44> 197 2150 385 c<94> p<35> p<34> p<32> p<38> p<43>
+ k<106> 383 p<24> p<67> p<27> p<33> p<39> p<31> p<37> p<46> p<50> p<25> p<53> p<59> p<26> p<45> p<57> p<69>
+ ICV_22 $T=0 0 0 0 $X=2540 $Y=356885
X2 VSS VDD 200 202 404 203 201 392 2180 254 391 2026 1600 2163 390 199 2164 2158 2029 205
+ 2028 2023 2192 419 2160 204 2193 2024 435 206 393 2162 2161 2039 255 394 2159 208 215 2165
+ 395 2169 253 207 399 209 2027 2166 2041 2040 2035 2059 228 412 2031 398 2175 2062 221 2167
+ 2032 2030 400 2081 218 2171 401 403 2043 2195 2170 402 2033 211 411 213 2174 2183 212 2034
+ 2037 2172 2036 231 405 1559 217 396 2046 442 406 214 1562 2191 2173 2025 2042 397 2182 2168
+ 224 2176 2045 407 409 210 408 2178 2044 220 1558 410 2181 219 2055 413 2185 2049 418 225
+ 216 2050 417 2177 2022 2057 433 2053 2052 1601 2212 222 227 223 2186 2047 2054 415 414 416
+ 2056 237 232 2179 2187 226 1560 2038 247 230 2189 422 2184 420 2063 2058 229 421 423 2060
+ 2051 233 2201 1564 235 234 444 2075 2061 236 251 2199 2196 239 2065 2194 424 429 426 2190
+ 238 427 2188 241 242 2070 436 2064 2198 425 454 1563 2048 428 2204 2200 244 2069 2197 2202
+ 245 430 246 2067 432 431 248 249 1561 2068 1602 258 441 437 243 438 2073 434 250 2071
+ 2066 252 440 2210 2074 2072 2080 2205 439 457 2206 2207 2076 2077 257 443 2203 445 2079 446
+ 263 256 459 261 447 259 240 2211 2083 448 2078 262 260 2082 2084 449 2093 450 451 2208
+ 2086 452 2213 271 461 453 264 2087 268 2214 455 467 266 265 2085 456 468 2088 267 458
+ 2217 462 269 481 270 460 2218 2222 464 463 2228 469 2227 474 2224 272 466 2226 482 2220
+ 2232 1961 495 2090 476 2215 2233 2229 1970 470 471 2231 2234 1566 472 473 475 2225 477 2216
+ 480 478 479 2235 2245 2153 1095 928 485 597 707 276 274 2155 275 112 483 484 1864 486
+ 2237 571 2239 2100 487 488 294 1565 491 2209 489 759 2246 2236 2097 2241 277 2247 2121 494
+ 128 278 279 493 497 290 288 340 496 295 492 498 2243 2242 1969 282 499 2240 500 501
+ 283 302 285 124 2223 502 2102 281 505 746 504 286 506 1046 528 2104 291 315 287 507
+ 512 378 289 508 509 510 490 329 704 2249 1074 122 513 514 2248 517 2251 293 2255 2252
+ 1044 2244 515 296 2127 531 511 520 518 304 2123 301 2107 2109 297 2115 344 1983 299 p<15>
+ 519 523 298 2250 1603 2253 524 522 p<7> 2221 153 2124 303 525 516 306 138 p<14> 157 2256
+ 305 376 526 503 307 308 530 309 333 310 k<78> 2230 2238 345 532 529 313 533 311 2263
+ 331 312 1987 2135 k<112> 534 609 2254 2219 p<8> 565 k<108> 348 172 332 140 2258 535 317 p<11>
+ 1991 314 k<94> 536 2140 316 539 538 594 545 1994 320 147 k<122> 2008 1647 540 k<115> k<91> p<27>
+ 541 p<24> 183 361 542 543 544 2142 p<12> 2261 2262 k<88> 2260 p<37> 330 547 549 550 321 1999
+ 323 156 551 1498 2259 1481 554 1077 552 322 328 557 566 327 1308 2004 324 325 1082 556
+ 555 326 2003 1604 p<26> 562 559 560 570 2147 166 563 564 1741 568 601 p<31> 2001 2006 k<95>
+ 558 567 2257 2264 p<16> 335 949 569 337 548 k<113> 572 339 346 343 341 356 336 342 k<120>
+ 573 k<46> 2266 576 k<107> 575 751 2146 577 2269 347 352 579 2267 580 k<109> 178 581 350 351
+ 1106 k<57> 355 583 2268 353 358 585 p<20> 587 582 584 2271 k<121> 591 k<101> 363 595 1092 359
+ 2012 2152 349 184 p<45> 596 k<89> 364 p<116> 2270 k<53> p<53> 600 588 p<25> 598 p<57> p<46> 599 771
+ 769 761 done 2156 2017 k<60> k<74> p<21> 605 k<28> 192 2019 k<114> 775 p<6> k<117> p<59> 610 379 553
+ 382 p<10> 381 k<116> 2272 602 1294 k<126> k<93> 608 159 2265 592 2020 p<23> 2021 384 k<61> k<103> k<100>
+ k<79> p<33> k<119> 383 k<123> p<5> p<18> k<118> p<2> k<104> k<105> k<124> k<127> p<0> p<13> p<19> p<9> k<106> k<125> p<3>
+ p<22> p<1> k<102> k<111> p<4> p<17> k<110>
+ ICV_24 $T=0 0 0 0 $X=2540 $Y=294165
X3 VSS VDD 390 616 391 2158 397 395 2168 409 2160 2159 617 619 2189 2165 393 394 406 618
+ 2161 2162 2179 392 2173 2166 2164 396 2163 416 398 621 2167 399 438 2279 2230 400 401 2175
+ 615 403 433 2174 2172 418 2171 404 405 620 2177 2180 2190 674 2182 408 411 2178 430 624
+ 2181 2169 2170 2184 410 2183 412 1601 441 1600 625 2176 413 626 414 643 2186 2187 2188 407
+ 2185 2273 417 415 2191 402 420 628 419 2196 422 631 632 2274 2194 423 443 2192 629 424
+ 421 2200 622 425 427 801 2198 634 2195 2193 2199 2197 638 428 635 429 2213 636 426 431
+ 639 2276 432 444 2203 434 1693 637 2202 435 2275 451 436 437 448 2206 641 642 2205 2214
+ 439 640 2201 2204 644 440 2277 2207 1602 445 1645 442 646 2219 648 2278 452 2210 447 2208
+ 652 455 651 450 449 2211 446 1968 650 2221 453 653 2212 2217 2098 655 454 654 2218 645
+ 623 457 2089 663 458 647 273 459 656 658 460 471 659 2284 2220 463 461 474 2095 462
+ 660 1967 2225 2222 2235 2094 464 2285 661 456 2224 473 466 662 2228 467 322 468 2227 470
+ 2226 477 2337 2286 849 2229 2231 664 469 1696 892 339 487 2295 2144 2232 2287 2288 2312 2282
+ 476 475 378 931 472 2289 2318 480 2233 478 2234 665 2296 481 2323 666 2292 2298 1092 2299
+ 482 1058 700 2290 479 488 1566 483 484 485 602 667 668 1020 2293 2280 2281 888 2096 671
+ 112 2104 1603 2291 670 495 490 672 2243 673 675 497 669 492 493 676 717 2297 1646 290
+ 491 679 288 496 682 677 678 507 2339 500 291 2101 284 680 684 2155 2250 1461 2300 504
+ 683 329 501 681 746 506 502 503 686 685 498 2099 691 2319 344 517 2313 526 315 687
+ 2108 505 2106 2105 2305 2249 2303 528 2087 688 508 509 690 510 2304 689 2302 511 692 512
+ 2306 2324 295 513 515 1045 530 523 2307 2310 516 1048 292 592 695 697 2247 2113 514 699
+ 518 2308 2309 522 694 550 553 953 2110 696 2301 520 2116 128 2111 698 1604 521 1981 2131
+ 701 k<87> 559 1982 703 2311 k<72> 713 705 k<73> 307 345 524 2254 2314 289 710 527 270 706
+ 533 2103 2315 708 2132 531 709 913 2316 1044 2093 1994 2125 711 2325 712 532 k<76> 573 2317
+ 2252 1647 722 2257 702 715 331 544 333 726 921 2136 2321 2129 2320 538 720 716 525 k<90>
+ 721 718 2322 719 144 2000 2261 693 1993 2259 725 2258 537 723 2130 558 542 724 541 539
+ 540 k<77> 2326 552 k<75> 729 2270 543 546 728 536 547 545 733 548 2327 732 730 293 731
+ 1996 549 560 551 555 2018 2264 575 736 734 321 2143 328 324 949 2329 1082 738 742 554
+ p<13> 561 556 330 557 564 2251 k<56> 382 190 2334 565 2331 741 563 740 935 2332 570 567
+ 1648 2007 2283 562 568 k<70> 361 569 743 183 744 338 745 2333 762 572 747 1741 k<67> 578
+ 2294 571 764 748 576 350 2268 1096 749 756 577 2335 950 581 727 2336 753 192 k<84> k<53>
+ 583 754 755 p<0> p<18> 580 752 2149 k<45> 579 582 k<69> 1480 k<64> 757 354 1111 587 758 k<102>
+ 759 k<68> 760 2004 591 360 k<82> 952 363 773 k<41> 761 593 735 k<74> 594 p<17> 595 2014 2330
+ done 597 p<50> p<39> 766 k<39> 596 765 186 767 2245 768 534 599 2338 k<96> 188 600 771 938
+ 374 k<57> k<71> 750 1120 p<4> 775 p<9> p<5> k<103> 774 195 304 310 k<63> 2341 k<98> p<19> 2340 776
+ 2342 365 2328 k<97> 2157 k<81> 610 714 k<80> k<65> k<62> k<55> k<54> p<2> k<85> k<83> k<59> k<78> c<78> k<93>
+ k<66> k<79> k<91> k<88> k<94> k<99> k<86> k<61> k<58> k<89> k<95> k<100> k<92> k<60>
+ ICV_28 $T=0 0 0 0 $X=2540 $Y=231445
X4 VSS VDD 780 818 617 781 782 628 406 2343 2344 793 988 2346 616 622 618 784 620 785
+ 790 619 809 2345 786 787 794 783 2353 789 2348 621 840 791 792 649 2354 2350 2380 2349
+ 803 990 795 630 635 796 625 633 801 816 797 2359 623 798 2373 2362 799 800 2355 810
+ 808 2352 624 802 2356 829 2357 2351 805 804 806 807 627 2358 2273 2347 817 626 2368 2360
+ 629 1693 812 1691 814 632 813 2361 631 2367 2275 2365 2366 815 819 831 822 820 825 634
+ 2363 823 824 788 2364 636 644 637 826 827 2276 828 1692 659 639 640 821 830 2371 2370
+ 643 2372 2369 642 839 2376 641 648 833 645 811 836 2375 2277 837 2278 2377 838 646 2374
+ 647 835 848 842 2378 845 650 843 651 2381 2379 653 652 844 846 465 847 2383 655 654
+ 2215 834 2382 656 1984 2092 658 2396 850 2384 851 684 852 2234 856 860 657 2398 2392 2223
+ 854 853 2385 858 857 1028 1030 859 2389 1019 861 2390 675 2388 867 1022 2391 663 869 664
+ 662 855 872 862 863 504 2387 666 864 877 865 2402 1014 1566 2395 868 870 1964 2393 1031
+ 2394 2403 871 2386 499 1025 880 873 2293 874 875 2291 668 879 667 866 2397 876 2236 2294
+ 878 2237 2239 1647 486 665 2399 2401 669 881 2240 2400 673 671 2241 2404 882 674 2242 307
+ 1694 493 494 2405 883 884 885 303 678 889 507 2244 291 756 886 528 315 290 746 679
+ 329 2303 2407 2248 2108 680 887 2406 681 683 682 677 890 891 892 931 893 685 2411 894
+ 686 895 896 1044 687 695 688 2305 689 2408 897 690 2111 898 2409 295 676 2300 899 514
+ 900 1048 692 901 2410 693 2414 2114 699 694 902 519 696 697 903 953 2429 714 2304 698
+ 2117 925 345 531 344 904 700 905 2311 701 702 703 906 907 2253 908 909 2412 1646 2121
+ 284 707 1286 704 2122 2313 529 2295 k<40> 706 910 2424 2126 2416 709 2310 911 710 135 2413
+ 766 708 711 2415 912 712 914 1695 k<34> 2328 915 133 916 2423 1391 k<37> 2418 2255 2417 917
+ 2320 716 918 2258 570 718 719 535 2249 922 920 1992 723 2420 2422 724 2421 725 2318 k<13>
+ 670 924 726 2154 2260 727 175 2425 926 728 2419 729 2327 927 112 2157 731 672 929 734
+ 2261 735 575 1696 2139 730 k<36> 933 k<49> 2141 913 k<66> 327 330 934 382 1697 k<39> 2427 2331
+ 936 738 740 940 555 939 749 741 288 324 742 744 322 941 745 321 743 943 357 747
+ 339 945 947 946 2333 944 343 2426 748 p<3> 581 948 k<67> 2267 1100 951 k<38> 179 754 2428
+ 753 k<7> 722 757 k<43> 585 1255 k<51> 2013 957 k<25> 760 759 568 713 762 done 2430 k<44> k<58>
+ 923 k<23> 2334 p<1> 565 956 768 c<95> k<24> k<48> 2151 k<42> k<21> 2245 360 769 600 k<45> 773 961
+ 605 k<31> 775 c<28> 962 2431 2272 601 k<59> 310 534 609 c<14> k<29> k<27> k<30> k<28> k<47> k<50> k<14>
+ k<41> k<35> k<32> k<33> k<46> k<52>
+ ICV_29 $T=0 0 0 0 $X=2540 $Y=200085
X5 VSS VDD 780 971 991 615 2347 2349 968 2432 782 786 784 2357 969 781 967 2343 622 785
+ 2369 783 979 2435 2434 2345 2346 982 787 788 2441 789 973 984 790 799 970 2436 2344 1692
+ 972 621 797 791 2356 976 792 800 818 2350 975 1691 1003 798 806 974 796 795 847 635
+ 2438 2352 2353 977 802 626 2437 804 801 840 985 2433 803 805 978 980 819 2358 981 807
+ 2378 808 809 823 810 811 986 813 629 1715 2351 2360 631 995 987 812 2364 846 990 814
+ 2365 826 815 1001 988 816 817 989 820 835 821 841 2363 824 822 827 2371 992 993 2377
+ 2366 994 2367 2275 2368 2439 825 2440 832 983 996 829 997 1693 833 998 2359 830 2419 999
+ 2354 2443 2372 1000 2442 2373 831 1002 1008 834 1004 2375 836 837 2446 2283 2376 1006 2444 839
+ 2445 838 1645 843 1007 842 2279 2379 1009 1010 845 2380 1012 1011 844 1005 873 2382 868 2381
+ 879 848 2450 850 1014 872 1013 1032 854 851 858 2391 853 2453 855 852 2386 859 1015 856
+ 860 2285 2447 1020 2389 1030 857 865 2388 2387 1016 1017 1022 1018 869 861 2448 1027 2396 867
+ 2449 1021 863 2397 2390 1019 862 2451 864 2395 2392 2452 2393 877 866 2399 1024 2394 870 1023
+ 871 1025 1026 875 874 2398 876 1028 1031 881 878 2401 1029 882 507 880 746 2454 506 557
+ 883 546 1034 1056 1033 884 303 344 2118 1035 677 1036 923 885 531 528 887 1037 315 1039
+ 2405 1043 1987 1041 1045 1040 1042 1038 715 898 890 1044 1047 1566 893 891 2307 1046 666 1048
+ 1049 894 897 899 1050 2306 295 1051 2112 896 1052 1053 900 695 903 902 1054 1055 2457 908
+ 2120 901 904 345 696 699 705 907 k<8> 2116 525 917 1057 2456 1059 909 2314 1985 1073 2458
+ 2455 k<9> 1986 910 1063 2105 911 2315 2459 1062 1064 287 135 1117 913 529 914 1066 k<15> 915
+ k<2> 2415 713 916 717 710 892 2096 1071 1068 1069 750 1070 919 2340 720 2460 922 1072 726
+ 2462 2138 1074 1058 2402 126 2461 k<36> 2265 2324 2463 112 924 1075 2466 2464 1991 938 2465 2148
+ 1076 554 1077 1697 1079 1078 731 2104 1084 730 2296 1080 2330 2262 1081 737 2467 1083 k<49> 932
+ 1085 2002 330 933 934 1086 382 936 2468 1109 935 937 1087 2469 1089 188 940 k<17> 1090 743
+ 2263 2261 941 943 k<35> 1093 1096 1091 1094 2005 2470 1095 928 k<38> 1097 945 946 2471 2429 2266
+ 574 944 1098 948 1099 332 2474 2472 1101 951 594 755 k<20> 1104 2473 1102 357 2299 k<18> 1108
+ 1107 2150 2290 2295 k<32> 1103 k<13> 1110 589 385 1113 952 931 k<10> 491 done 1111 2271 k<25> 953
+ 1114 k<0> k<33> 2475 1115 c<124> 2404 598 956 2478 2476 2477 764 371 771 2479 k<16> 566 2335 2133
+ c<117> c<121> c<127> c<125> 1123 k<26> 327 608 1124 k<22> k<3> k<21> k<6> k<12> k<4> k<7> k<19> k<27> k<11> k<23>
+ k<14> k<24> k<5>
+ ICV_30 $T=0 0 0 0 $X=2540 $Y=168700
X6 VSS VDD 2280 1009 2507 1318 1130 2209 2484 967 1128 2216 1133 2480 1137 2518 2483 2482 1129 968
+ 1962 2485 2502 969 1006 2351 2481 1131 2348 1134 1729 625 1132 1149 2497 2498 1136 2501 1135 2492
+ 2490 1139 2493 2281 1140 1138 2496 989 2400 970 2519 2499 2489 2488 1322 2500 973 2516 1141 2494
+ 794 2503 1142 2486 2505 2487 2432 1143 2509 972 1146 1145 2520 2495 2504 792 831 1732 2273 2511
+ 1144 2508 971 1147 2510 974 2542 975 2513 1148 1159 816 2434 1325 1000 1731 2521 780 2514 1150
+ 2540 2444 2433 2361 2541 801 2442 812 977 2515 2517 2528 2525 2512 2355 976 1336 978 621 1152
+ 1151 2491 1153 979 2527 2506 983 2524 2536 980 1161 1154 2544 1155 2522 1156 2526 2529 2523 1157
+ 643 1158 981 2531 2354 2360 2534 2530 2435 1162 2532 2367 982 1165 2535 2533 1692 986 2440 808
+ 1163 2537 1004 1164 1975 2362 631 2539 2436 2538 2543 987 1166 1167 984 2428 2275 1168 1169 988
+ 2545 1007 2374 1170 1160 2546 1171 2437 2547 1172 990 2359 1973 1173 2466 2438 2274 992 622 2556
+ 110 1176 995 2552 993 1177 2554 1374 994 2570 2553 1733 2551 2555 786 2603 1002 2558 2557 2565
+ 998 1977 1179 2370 1187 1180 828 2580 991 2439 1174 1181 1182 1375 997 2559 999 2446 2562 1186
+ 996 2419 1185 1978 1184 1183 2561 2573 2563 2589 1378 1001 2569 2564 2568 1003 2567 1734 1178 2560
+ 2572 2571 1189 2550 1188 2575 2443 2548 1190 2445 1005 2441 2283 2574 1191 1199 2576 2566 2578 2581
+ 2595 2577 2582 2587 1192 1008 1193 1735 1175 2584 2585 2549 1194 2282 1736 2586 2583 2592 1011 1010
+ 1195 1196 1197 2590 1377 2579 1737 1012 1198 2591 1202 2594 1972 1976 849 2593 2384 2604 1200 2602
+ 1209 476 2588 2597 1201 2385 1203 1014 1206 2596 2383 2091 1204 2598 1205 858 868 2599 1013 2284
+ 1022 1207 661 1015 854 1208 2600 660 473 872 1030 2452 869 1018 1964 1016 2447 2601 2453 1017
+ 1211 1019 1212 1210 2387 2449 2448 861 1566 2608 2450 1214 1213 2465 2389 1215 1216 1225 2287 855
+ 1020 666 2607 1218 2390 2451 2393 879 1027 1224 1220 1021 1221 1222 2232 1023 2288 1219 877 2244
+ 746 1243 1223 1226 1024 472 2626 480 1227 1237 2238 2610 1028 1025 1026 874 2398 2289 1229 1231
+ 1258 1230 2611 2292 1238 1228 1233 1029 1031 2297 1032 2401 2399 1738 873 2621 1101 1234 1235 2612
+ 1236 2615 2613 1249 1239 546 2454 1463 1240 1241 2403 1054 2614 731 303 1034 1242 1472 2298 2617
+ 1035 1299 1244 2605 1248 1037 1245 1036 2616 507 1246 1247 714 1048 2455 288 531 2301 1041 295
+ 2620 528 1038 329 315 888 1250 1039 1251 2618 1040 2409 715 2117 1033 1043 2302 890 1044 895
+ 2407 1042 1051 1045 691 695 1047 2622 1046 1257 2619 1049 2408 1252 1050 2456 147 1253 1254 1052
+ 1053 1269 513 2457 1266 1303 1256 698 1259 905 925 1260 1057 1261 1262 906 1058 2114 1061 1263
+ 1988 2318 345 2340 1056 913 914 1273 2312 1264 k<2> 911 k<9> 284 1265 1062 2623 1267 2256 1064
+ 909 912 711 k<1> c<104> 1268 1272 2316 2624 2317 1066 1255 1271 1063 2625 2417 1270 917 287 1864
+ 1274 2322 1275 k<12> 720 920 1069 2249 1276 921 k<5> 1465 1277 1995 2323 670 1279 1281 1280 1072
+ 1068 1073 1278 721 112 c<119> 1282 696 2423 1075 2246 c<108> 699 2628 2627 k<11> 1284 1390 175 1283
+ 2020 1285 926 1084 726 2631 2134 730 1286 732 1287 1076 1077 1078 1288 1289 733 2630 1079 710
+ 2330 2629 736 2632 1290 562 1081 1085 k<17> 1080 773 1291 1292 1087 2329 1294 583 k<20> 1088 1083
+ 1293 557 k<32> 1740 1297 554 1301 1086 c<122> k<52> 2633 188 588 584 1089 349 1090 2634 1091 2011
+ 941 1295 1092 2326 1296 745 k<4> 2635 1298 1106 1093 580 944 2472 943 2017 1096 2638 1097 1307
+ 1104 1302 1098 761 751 928 1739 1103 949 k<50> 1304 2636 1102 2270 k<38> 2637 2015 950 901 1310
+ 2295 357 722 1305 2473 2467 1109 1311 940 c<112> c<123> c<103> 1110 2639 2640 1306 2104 2471 k<3> c<102>
+ 939 c<96> 1113 765 2327 2464 2096 c<115> 1114 c<100> c<99> 942 c<109> c<101> c<126> c<114> 300 2641 c<111> c<98>
+ 671 done c<118> 2430 c<97> 1309 c<113> 1074 c<90> 569 c<120> 2105 2004 c<83> 774 2338 1120 2642 1312 c<107>
+ c<84> c<116> 2468 c<110> c<89> k<19> c<87> 1123 c<105> 776 c<106> c<88> 2341 2431 c<91> c<85> c<77> k<0> 1124 c<82>
+ c<30>
+ ICV_32 $T=0 0 0 0 $X=2540 $Y=106005
X7 VSS VDD 1324 1321 1316 2480 1315 1130 2645 2502 1332 2482 1129 2510 2483 2663 1318 1149 1317 1131
+ 1128 2490 2484 2489 2495 1135 2485 1729 2487 1139 1142 1132 1337 2491 2488 1326 1133 1731 1134 2644
+ 2494 2643 2505 1145 1320 2508 1322 1136 1138 1323 2493 2652 1331 2499 1140 2512 2492 2496 2498 2507
+ 1141 2500 2646 2648 2653 2659 2649 2647 2497 1147 1319 2504 1329 1143 2501 1144 1137 2651 1338 1327
+ 1146 2654 1325 2656 2506 2655 2509 2660 2513 1349 2521 2511 1157 1730 2650 1328 2662 2514 1161 2516
+ 2517 2400 2668 1334 2661 1150 1330 2657 2535 1348 2518 1335 1151 1156 2520 1347 1340 2658 1333 1153
+ 2536 2525 2522 1339 2523 1336 1152 2524 2519 2530 1148 2666 2527 2664 1166 2533 1159 1155 2531 2528
+ 1158 1341 1346 1344 1160 2526 2534 1342 2529 1343 1162 2532 1345 2665 1163 1164 1168 2540 2537 1732
+ 2669 2539 2667 1167 2541 1352 1350 2538 1165 2670 1351 1169 2546 1170 1353 1154 1357 2544 1361 1354
+ 1365 1369 2561 1174 1364 1172 1356 2551 2550 2548 1359 1175 1179 1358 2554 1185 1176 1362 2555 1363
+ 2598 1360 1177 2671 1355 2672 2553 2552 2559 2673 2577 1370 2675 1784 1178 1733 1375 1783 2557 1368
+ 2674 2556 2677 1182 2564 2569 1181 1180 1210 2579 1204 2558 2568 2678 2562 1183 2676 2560 2571 1184
+ 2684 2563 1189 1366 2681 1367 1186 1373 2566 1734 2565 1192 1187 1202 1188 2567 2547 1190 2570 2572
+ 2573 2578 2576 1379 2575 2574 2680 1193 2679 1371 1191 2581 2580 2688 1374 2582 2593 2588 1173 1198
+ 1735 2682 2683 2584 2583 2587 1194 2589 1195 1196 2590 2586 1736 1372 1376 2591 1211 1197 2685 1387
+ 1199 2592 2691 1380 1200 2599 2594 2687 1378 1201 1203 1383 2596 2689 1205 2595 1382 1381 2686 2690
+ 2597 1388 1206 1208 2601 1207 2693 2600 2692 1384 1385 2606 1390 2605 1209 1389 2602 2603 1386 1391
+ 2694 2604 1212 1213 1214 1392 1215 2695 1216 1394 2696 2609 1393 1218 2707 1419 2286 1217 1395 1401
+ 1396 2698 1219 1397 2699 1398 2697 2612 2608 1220 1222 1409 1223 1221 2610 2700 1235 1400 1405 1399
+ 1408 1226 1411 1225 1785 1402 1228 1227 1403 2701 2711 1230 1404 1239 1224 1229 2706 1406 2705 2704
+ 1232 2611 2703 2702 1233 1247 1231 1426 2720 1236 2708 1407 2709 1410 1416 2710 1240 2613 1425 2712
+ 1413 1422 1412 1234 1414 1245 1415 2713 1237 2715 1446 1238 1417 1418 2719 2738 2714 2725 1420 1241
+ 2717 2718 1421 1248 1424 2716 2734 2614 2721 1430 1243 1244 2722 2615 2724 2723 2616 1427 1423 2727
+ 1428 1429 1434 1431 2730 1246 2726 1242 1249 1432 1250 1786 1440 1433 1435 2618 2729 2728 2617 1436
+ 1441 1251 2732 1439 1437 1438 2731 691 1442 1252 1455 2620 1456 1447 2733 1443 1444 1445 2735 1255
+ 1448 1253 1453 1254 1459 2736 1450 315 2406 1449 1256 1258 2410 1451 2411 1739 1257 2737 1260 1259
+ 1458 905 1452 1261 1460 2412 1454 1263 2458 1051 1265 c<73> 1048 1264 1457 1262 2465 1271 1266 1303
+ 2459 2413 1461 1269 1268 c<65> 2623 1462 c<66> 2319 916 1267 1275 1280 1695 2417 1273 1274 1464 918
+ 1276 528 2416 2418 1463 1279 c<69> 1070 c<72> 2626 1469 718 1277 1278 2128 1281 896 2461 1071 2422
+ c<76> 1283 1466 2462 1285 345 1467 1284 2464 1468 1035 2635 1286 1287 2425 157 1696 1044 2622 2424
+ 2621 1289 k<6> 531 1290 2630 k<4> 1306 1056 2009 1471 1037 1472 1095 1740 2739 1470 1293 2632 1291
+ k<3> 2631 1473 2290 1294 1292 1741 1475 2426 2634 1474 775 329 2469 2333 2471 1295 1297 1296 1487
+ 1300 1481 1299 1476 1298 1477 1094 2740 1301 751 1302 947 1111 1478 2637 1304 2636 1479 489 752
+ 1101 1482 1100 2337 2325 k<18> 1106 722 1490 2414 1305 c<43> c<44> 2479 2145 1485 c<38> 2638 c<62> 758
+ 1483 1082 c<35> c<54> done 2474 1307 c<58> 2619 2119 2329 358 1308 2137 2269 1099 2308 571 2336 c<42>
+ c<50> c<46> c<47> c<60> c<32> c<49> c<33> 1117 c<80> c<40> c<57> c<52> c<59> c<75> c<61> 1309 c<56> 1310 c<70> 2478
+ 2309 c<67> c<51> 2339 1115 1311 2463 c<63> 1648 c<31> 1104 c<81> 1492 1312 c<39> 1493 962 c<71> c<48> c<68>
+ c<55> c<41> 2342 c<53> 2477 c<74> c<45> c<64> c<29>
+ ICV_35 $T=0 0 0 0 $X=2540 $Y=47100
X8 VSS VDD 2481 1315 1317 2490 1316 1133 2660 2486 2484 2653 1129 1319 1330 1324 2487 2643 2498 2494
+ 1321 1320 2644 2655 2646 1318 1128 2650 2658 2502 1323 2661 2645 1337 2648 2509 1328 1148 2503 2647
+ 1322 2664 2659 1144 2656 2515 2489 1325 2649 1339 1326 1349 2511 2652 2654 2651 1327 1329 2535 1335
+ 1131 2657 1341 1331 1340 2668 1332 1333 1334 1350 1336 1154 1347 1130 1338 1159 2534 2662 2507 1344
+ 1342 1343 2665 2663 1352 1345 1346 2667 1353 2666 1348 2670 2669 2552 1351 2543 2542 2545 1360 1171
+ 2693 2547 1355 1358 1356 2549 2682 1354 2673 2686 1361 1363 1362 2671 2674 1783 1375 2675 1357 2684
+ 2569 1784 2677 1364 2571 1190 2676 1380 2570 2678 1365 1386 1367 2687 2566 2672 1368 1734 1376 1359
+ 1389 1184 1369 1370 1383 1195 2680 1371 2679 1366 2681 1372 2580 1373 2683 2694 1379 2585 2685 1374
+ 1737 1377 1378 1382 2605 1381 2690 2688 2691 2606 2689 1384 2692 1385 1388 1387 1390 1391 1393 1392
+ 2695 1394 1396 2733 2607 1397 1395 2697 2698 1402 2696 2702 2617 1404 2700 2710 1403 1398 2699 1399
+ 1401 2701 2722 2705 1405 1412 2704 1444 2703 1406 1407 2706 2712 2707 2709 1416 1411 2716 1408 1413
+ 2714 2713 1410 1414 1425 2715 2737 1236 1415 2730 2719 2711 1418 1417 2717 1217 1420 1438 2718 2721
+ 2728 1421 2720 1422 1429 1423 1424 1426 1433 2723 1427 2724 2726 1430 2708 1431 1435 2725 1432 1441
+ 1428 2620 2609 1785 1437 2727 2731 2729 1455 1453 1436 2732 1439 1449 1445 1400 1442 1448 1450 1443
+ 1419 2736 2735 1786 1446 1447 2616 2734 1434 1452 1451 1454 1459 2738 1440 1457 1458 1456 1460 1462
+ c<15> 1272 1270 1059 2625 c<8> 1463 1464 c<1> 2624 1465 c<12> 2321 c<2> c<9> 2460 1466 2465 2420 c<16>
+ 1461 1266 1282 2421 c<5> 1468 1467 2627 c<11> 2629 1469 2319 929 1288 1477 1291 1470 1472 2739 1478
+ 1473 1051 1474 1303 1476 1265 1475 2332 2470 1480 c<24> 1099 957 2633 1479 1481 1482 1107 c<17> 1108
+ 1106 1483 c<34> c<36> 1471 1485 c<4> 2740 c<6> c<37> 1487 c<3> 2641 c<10> 1490 c<25> c<18> 2639 2475 c<20>
+ c<23> 2427 2640 c<7> c<13> 961 c<22> 2628 c<19> 1492 1493 c<26> c<21> 2642 2476 c<0> c<27>
+ ICV_36 $T=0 0 0 0 $X=2540 $Y=210
.ENDS
***************************************
